<svg:svg xmlns:xlink="http://www.w3.org/1999/xlink" xmlns:svg="http://www.w3.org/2000/svg" version="1.1" width="595px" height="842px" viewBox="0 0 595 842"><svg:g transform="matrix(1 0 0 -1 0 842)"><svg:defs ><svg:style type="text/css">@font-face { font-family: &quot;g_font_3&quot;; src: url(data:font/opentype;base64,AAEAAAANAIAAAwBQT1MvMmLSWIkAAADcAAAATmNtYXDCjyO8AAABLAAAAIRjdnQg+z6j2gAAAbAAAAdaZnBnbQjouigAAAkMAAAF12dseWYQL03UAAAO5AAAQ5poZWFk58I9qgAAUoAAAAA2aGhlYRJ+FiYAAFK4AAAAJGhtdHhZvsAMAABS3AAANXRsb2NhA3h0DgAAiFAAADV4bWF4cBVHAbMAAL3IAAAAIG5hbWX+r+oRAAC96AAAAmpwb3N0AAMAAAAAwFQAAAAgcHJlcPFK5RYAAMB0AAAR0gAABAABkAAFAAAEAAQAAAAEAAQABAAAAAQAAGYCEgAAAQEBAQEBAQEBAQAAAAAAAAAAAAAAAAAAAAA/Pz8/AEAAIAB5CAACAADMCCQEAgAAAAAAAQADAAEAAAAMAAQAeAAAABoAEAADAAoAIAApADkASQBQAFUAWQBbAGkAcAB54AD//wAAACAAKAAuAEEASwBSAFkAWwBhAGwAcuAA////4//j/+P/4//j/+P/4//j/+P/4//jIAMAAQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABboAHAW6ABwFpwAcBCYAHAAA/+QAAP/kAAD/5P5p/+QFugAc/mn/5ALqAAABHQAAAR0AAAAAAAAAAACyAKwA1wEoASAAswH6ABcA+AEZATEASQAEAPcAAwCvAP0AlQAUAFQAlgESACQAFgBVAEkBBAEZASsAjAGb/3b/6QA9AJIAov+3AYL/qgAWAI8AxgD4ABwA3gQBADcATgBVAFUAZQDpA+UAWf+aAAgAhwALADsAUgEWAGEA1gDWAPUAAACTAJQAvgF8//gABAAUAIIAkgA8AEEAQf/B//wAKgCMBJAF2Am1AJEAuwEG/2P/aQAeACIAigIr/9b/3wAmAFkAowCsAQQBKwHABEgAIQBrAIUAmAEZA8YAawCVAKQA/gEMAl0DQwW/AAAASQBWAG4AdwCKAKoAygESAVAF2AXw/3v/5wAGABMAKABhAGkA6QE1AU0CpQQM/z7/2gBbALkAyAEZARkBGQHABFsEpwVb/j//nf/CABUAtwEKAbwBwQUyBY79gf+h/64ADAAmADEAPQBOAFYAYgCDAMEAyQDxAPICf/9/AEgAUwB3AMUBHQEgASYBKAHWAhkCfgJ+A9MALgBBAF0AawB1AJ8AsACyALoAuwC9ANYA2wDgAOUBFAEbAUoBYgGRAfICDAJkAs8DmwO0A9QEAQSpABYAIwAlACoAdAClALYAzADNAM8BBQEgATABUAFqAW8BlwGdAeACsALsAvcECASDBPsE/QUm/uD++/9O//UAGAAaAEwAegB/AJEAowCzALQAzgDVAPIA8wD2ARABOAFoAaEBsAHgAewCCQIiAk8CcAKWAqUCrQNOA5EDwQQ1BEIEawTNBNoFhgWLB2EH/vym/pP+rf7R/7f/0QADAA4AGAAmAEYAaQCBAI8ApQC/ANMA1QDZAN0A4gEZASsBOAE7AVoBXgFoAXMBiAGUAa0BxQHRAeoB8gIAAgACAAIiAjsCRAJPAm8CcgJ+AoICkwKUAqUCzwLPAtAC2gLdAusC9QMFAyIDNgNxA6EDsAO4A9AD5gQQBCYELgQxBE8EWgT/BTIFMgVHBVMFqAWrBcIF8AY8BmQGcAboB4IHhAjM/Sr93v4A/mj+sP6z/6oACABZAHoAkQCeAKIArwC0ALsAygDMAM4A2QDgAPQBFAEaASEBJwErATkBRgFLAU0BVwFcAWUBggGHAZIBmAGbAaIBrgHFAcUB0QIHAiICKwJBAlMCYQJlAoQChwKNArQCtAK6AskC1gLYAu0C9QMXAyMDKwMxA0kDWgNbA24DcQN0A34DhAORA5EDqgPPA9MD5wPoA+0ECAQXBB4EdQR6BJkEpwS0BNEFTAVtBW0FogW/BcAF0QX8BfwGAgYaBhwGLwZqBqgG4gcGBzYHUAeJB9QH8whwARwBKgEaASAAAAAAAAAAAAAAAAACGQALAB4CqgIUBH8B7QAAAB0BBAAPAJEAKwGIAVMBEgHzAD8D/gFoAQ4EfwHtA24DFQIZBBMAAAAABkAEsAAAAnQBuwA1AcUAfwYCAwEAAATgALIB3ALgBMMCPQDVAWABGQSnA24FygIhAKsEJgCQArwCuwFCALQCPAJWApwDAAHlAagA5QBrAHgAlAFrAXMAqwHtAToBfQE3AX8A1AIWA1MBhAA8/6ICBAEJAUkB8ABuAxUAgQRkAF4AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABOQDcAOn+ngQNBHwBKwC4AJYAWQCsAN8BqQD6AQX/7AAXAAMAVQBhAAQAjACjAIUAKAEgAF0A1gB/ASYBGQEEAWwGzwC0AQYAAAc3Bj4EegDwAPkA6QW6BCYEQgAA/+f+aQSeBOP/N/8tASABBQEgAKgAdABoAEcA8gDlANkAvQCoAGgARwBcAEgACgAoADIAQQBQAFoAZAB9AIcAkf+w/5z/g/95/28AywEgAPoBLAH6AaAA1QC4AFwAPADIAMgAjwDZAYsAswBHAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA/mQAwADqARgBJQEyA7AD7QV2BZAFqgW0Bb4FzQYxAHgAhACbAMwA4gD0AQoBIAFjANEA6gD3AQgBQgAZACwANABBADgASABYAGwCWQO9AEMBGgBwANMAKAA3AEIAUABaAGQAcwB4AIIAjACcAKUAvQDOAPABEAFcAL4A2AECARcBLAFjAOoBCABBAEsAVQBfAHMApgEJAYMBswBBAGQAHgAqAOsA+gEOATgCdAAsAEAAggCWALYAwADMANwA5gDwAP8BCgEgASwBOwFEAVYBYwD3AFcAZAEQATYAUAGxAAD/tgA5AE4ARAPMAOUAJAEQAEIBIgGkAPAAYADgAA4AHQA5BeMBAgAs/k7/OAJpA70BFgD/AA4AoABUABsAPQFxAEEADwBQAP0AFQFPADX+UgAsANMBAwSwAdIAtgDAAJkCZf+HA3f+bADLAKkAXABABHYHRAAAQEFUQD8+PTw7Ojk4NzU0MzIxMC8uLSwrKikoJyYlJCMiISAfHh0cGxoZGBcWFRQTEhEQDw4NDAsKCQgHBgUEAwIBACxFI0ZgILAmYLAEJiNISC0sRSNGI2EgsCZhsAQmI0hILSxFI0ZgsCBhILBGYLAEJiNISC0sRSNGI2GwIGAgsCZhsCBhsAQmI0hILSxFI0ZgsEBhILBmYLAEJiNISC0sRSNGI2GwQGAgsCZhsEBhsAQmI0hILSwBECA8ADwtLCBFIyCwzUQjILgBWlFYIyCwjUQjWSCw7VFYIyCwTUQjWSCwkFFYIyCwDUQjWSEhLSwgIEUYaEQgsAFgIEWwRnZoikVgRC0sAbELCkMjQ2UKLSwAsQoLQyNDCy0sALAXI3CxARc+AbAXI3CxAhdFOrECAAgNLSxFsBojREWwGSNELSwgRbADJUVhZLBQUVhFRBshIVktLLABQ2MjYrAAI0KwDystLCBFsABDYEQtLAGwBkOwB0NlCi0sIGmwQGGwAIsgsSzAioy4EABiYCsMZCNkYVxYsANhWS0sRbARK7AXI0SwF3rkGC0sRbARK7AXI0QtLLASQ1iHRbARK7AXI0SwF3rkGwOKRRhpILAXI0SKiocgsMBRWLARK7AXI0SwF3rkGyGwF3rkWVkYLSwtLLACJUZgikawQGGMSC0sS1MgXFiwAoVZWLABhVktLCCwAyVFsBkjREWwGiNERWUjRSCwAyVgaiCwCSNCI2iKamBhILAairAAUnkhshoaQLn/4AAaRSCKVFgjIbA/GyNZYUQcsRQAilJ5sxlAIBlFIIpUWCMhsD8bI1lhRC0ssRARQyNDCy0ssQ4PQyNDCy0ssQwNQyNDCy0ssQwNQyNDZQstLLEOD0MjQ2ULLSyxEBFDI0NlCy0sS1JYRUQbISFZLSwBILADJSNJsEBgsCBjILAAUlgjsAIlOCOwAiVlOACKYzgbISEhISFZAS0sS7BkUVhFabAJQ2CKEDobISEhWS0sAbAFJRAjIIr1ALABYCPt7C0sAbAFJRAjIIr1ALABYSPt7C0sAbAGJRD1AO3sLSwgsAFgARAgPAA8LSwgsAFhARAgPAA8LSywKyuwKiotLACwB0OwBkMLLSw+sCoqLSw1LSx2uAI2I3AQILgCNkUgsABQWLABYVk6LxgtLCEhDGQjZIu4QABiLSwhsIBRWAxkI2SLuCAAYhuyAEAvK1mwAmAtLCGwwFFYDGQjZIu4FVViG7IAgC8rWbACYC0sDGQjZIu4QABiYCMhLSy0AAEAAAAVsAgmsAgmsAgmsAgmDxAWE0VoOrABFi0stAABAAAAFbAIJrAIJrAIJrAIJg8QFhNFaGU6sAEWLSxLUyNLUVpYIEWKYEQbISFZLSxLVFggRYpgRBshIVktLEtTI0tRWlg4GyEhWS0sS1RYOBshIVktLLATQ1gDGwJZLSywE0NYAhsDWS0sS1SwEkNcWlg4GyEhWS0ssBJDXFgMsAQlsAQlBgxkI2RhZLADUViwBCWwBCUBIEawEGBIIEawEGBIWQohIRshIVktLLASQ1xYDLAEJbAEJQYMZCNkYWS4BwhRWLAEJbAEJQEgRrj/8GBIIEa4//BgSFkKISEbISFZLSxLUyNLUVpYsDorGyEhWS0sS1MjS1FaWLA7KxshIVktLEtTI0tRWrASQ1xaWDgbISFZLSwMigNLVLAEJgJLVFqKigqwEkNcWlg4GyEhWS0sRiNGYIqKRiMgRopgimG4/4BiIyAQI4q5AqcCp4pwRWAgsABQWLABYbj/uosbsEaMWbAQYGgBOi0ssQIAQrEjAYhRsUABiFNaWLkQAAAgiFRYsgIBAkNgQlmxJAGIUVi5IAAAQIhUWLICAgJDYEJZsSQBiFRYsgIgAkNgQgBLAUtSWLICCAJDYEJZG7lAAACAiFRYsgIEAkNgQlm5QAAAgGO4AQCIVFiyAggCQ2BCWblAAAEAY7gCAIhUWLICEAJDYEJZWVlZLQAAAgEAAAAFAAUAAAMABwBCtAIB/gYHuAI/QBMABQT+AwAKBwT+AQAZCAYF/gIDvAEmAAkBsAEYABgrEPY8/TxOEPQ8Tf08AD88/TwQ/Dz9PDEwIREhESUhESEBAAQA/CADwPxABQD7ACAEwAAAAQBr/lECaAXTABAARkAOKA+nAwIICQEACRAAEgi9ASIACQABASIAAAKUQAoJ8wybIAQwBAIEuAKWsxGlaxgrEPZd7f307RDtAD8/EDwQPDEwAV0BIyYCNRATNjczAgIVFBIXFgJlwZmgY1aEwIlnPTUj/lHnAfLpASEBAuC9/tH+V+6k/qibZgAAAQBD/lECQAXTABAASUAYJwInCmcCZwqXAqcCqA4HCQgQAAgQABIQvQEiAAAACQEiAAAClLQI8wWbDLgClrMSakMYKxD27f3k7RDtAD8/EDwQPDEwAV0TPgM1NAIDMxYSFRQHAgNFU0Q6HGaJv5enQkus/lGyvvjfde4BqQEv1/4e+NHv/vT++wAAAQCTAAABrAEZAAMAJEAVAjgACgImDwAfACAAMAAEABkEZ3YYK04Q9F1N/QA/Te0xMDMRIRGTARkBGf7nAAAB//3/5wI7BdMAAwA4QB0AAQFJAgMUAgIDAgEAAwAKAesCGgUD6wAZBJNsGCtOEPRN7U4Q9k3tAD88PzyHBS4rfRDEMTAHATMBAwFr0/6RGQXs+hQAAAIAVv/nBA4FwAAOACAAk0BLeAqICqcBqgeqCacOtwnICQhWEVkWWRpWH2cRaBZoGmcfCDkCOQY2CTYNSQJJBkUJRg2nCcsCyQbECcQN2QLbBtQJ1A0REBggGAIYuP/AQCUSFjQYpggNHw8vDwIPQBIWNA+mAAUd2E8EAQQaIhTYCxkh08IYK04Q9E3tThD2cU3tAD/tK3E/7StxMTABXQBdXQEyFxYREAcGIyIAERA3NhciBgcGERAWFjMyNjc2ERAmJgIy1XiPkHfV1v76kHfVM1AWHTRPMzNQFh00TwXAmLT+X/5gtpYBSQGmAZ62lulBVG3+/v7+wUBBVGwBAgECwUEAAQCiAAADJgXAAAkAVkAJawJ7AosCAwIEuAEps18FAQW4Al63CAkFAQAMCQC7AVgAAgABAl1ADQUABB8EIASwBAQEGQq6AacBoAAYK04Q9F08TfY8/TwAPzw/PPRd7TkxMABdISERBgc1NiQ3MwMm/uea0W4BAjDkBCOQRf8kyYYAAAEAMwAABAwFwAAdAT9AX7UYthq5G8oExxjQGNAZ0BoIQxtDHEMdVhmbBJUYqgSmHAgGGiAAKAY3GkgEQxhDGUMaCCQYJBkkGgMWJgRWBIgYnBucHJwdqhyqHQgSAB0QHSAdMR12HYQdkB3WHQgduP/AQBYUFTQdAhAMDx0QACAAAiAAMABAAAMAuP/AsxIWNAC4AqGzAgEMD7gBVkAjHwwvDAIMQBIWNAymEwUJ2BYWAU8AAQAaHw/YEHcCGR7TwhgrThD0TfTtThD2cTw8TRDtAD/9K3HkPzz9K11xPBESOQERMytdQ1xYuQAd/8CyETkduP/Asg85Hbj/wEAOEDkECBA5BQgROQQIETkrKysrKytZsQYCQ1RYQAsJGxkbAhsTAQQTAAAREjkREjldWTEwAV1LUVi9ABv/4AAc/+AAHf/gODg4WQFxXV1dAREhNhI3Njc2NTQmIyIGByU2JDMyFhUUBgcGBAYHBAz8JxCg7L4rOmVZWGgI/ugZAQjG2fhHTTP+9kcWAQX++5QBCduxP1dVXmVqexzoyuquY7NiQfRQJgAAAQBN/+cEGwXAACkA2UAyhxXJFQJ7HIscAqYDqQWnFLYDugW2FNoY3RkIFhQBjRaNFwIhCg0ABAEXExYhHw0QDAq4ASRADE8NAUANjw0CDQ0BFrgBAkAPHxMvEwITQBIWNBOmGwUBuAFWtRAEIAQCBLj/wEAyEhY0BKYnDbAMwAwCDAwWENh/H48fnx+vH78fBR/gB9hPJAEkGisW2Bd3AdgAGSrTwhgrThD0Te307U4Q9nFN7fRd7RE5L10AP/0rceQ//Stx5BE5L11x7QEREjkROQAREjkREjkREjldMTABcV1dAF0TJRYWMzI2NTQmIyIHNxY2NTQmIyIGByU+AjMyFxYVFAcWFhUUACMiJE0BEA1yUVd3clI2Sx9yeFhJSGYL/v0bbcN5z31n036X/ubSx/76AYUhaG6EcGp8FeUDaVdKWGRgLIWfW4RsiMFzG7yFwf7w5QACACYAAAREBcAACgANAN9AOQwgDTkJDBkMKwxTDGsM4gwG7Q0BBgQWBCUEKA1IDVsNpw23DcYNCQECCAAMBg0HBQoLDQcADAwNDbgBrkAaAwQUAwMEAwIMBA0DDQIECgAHQA3ADdANAw27ASgACAACAbS2AAQEAAwMALgBWLQFjwoBCrgBAkASEAefB78HAwcaDz8CfwICAhkOugFMAUgAGCtOEORxEPZdTfRdPP08AD8/EPQ8/V08ARESORI5OQAREjkSOYcFLisEfRDEDw8PsQYCQ1RYQAstDD0MTQzNDN0MBQBdWTEwAV1dAF0rIREhNQEzETMVIxEBEQECfv2oAnzstrb+8P6vASf2A6P8Xvf+2QIeAfX+CwABAFv/5wQ1BaYAHQEQQCkIDiAMNxJFEkkZmQ2eDpcS2g4JEhETEiERIxKFEgUABAENCgwMDRIREbgCoEAWDg0UDg4NEgoUIAEwAUABA1ABkAECAbgBVrUQBCAEAgS4/8C3EhY0BKYbDQy4AlpADR8KLwoCCkASFjQKphS4/8BACxQWNCAUMBRAFAMUuAGrQBQRER8QLxACLxA/EE8QAxBAEhY0ELgCoEATDw8OBA8Q4AfY0BcBQBcBFxofDrgBIUASDXcBvNAAAUAAnwCvAAMAGR7TuQFHABgrThD0XXFN7fTkThD2XXFN7fQ8AD88EP0rXXE8EPZdK/0rceQ//Stx5F1xERI5hwUuKw59EMQBETkAERI5ERI5MTABcV0TJRYWMzI2NTQmIyIHJxMhESEHNjMyABUUBwYjIiRbARgMdk1YenlheWDkkALn/e4sXmK7AQRpj/7L/wABeR1fb4+Qh4drIQL7/vn5L/7w2bWOwtoAAgBX/+cEKgXAABcAIwC9QDtqC3UIhwiXGacFpwipDqoTuQ62Eb0TwBHPEw0VBTYRRBB6FrUC0hDQFAe7AM8AAgAEAQcYEhAbIBsCG7j/wEAeEhY0G6YPDR8hLyECIUASFjQhpj8JAUAJ0An/CQMJuAFPs68BAQG4ASFAIh8ELwQCBEASFjQEphUFAdgAdx7YTwwBDBolGNgSGSTTwhgrThD0Te1OEPZxTe307QA//Stx9F32XXHtK3E/7StxARESOQAREjldMTABXQBdAQUmJiMiBgc2MzISFRQAIyIAERAAMzIWARQWMzI2NTQmIyIGBA/+8ApUQ1l7EGmcsPv++M/e/uIBKu6n2/2hflFOaHBUUXAEUx5UUKD9fP701OH+8AFZAYkBkwFku/zpiZV6i4+FfwABAFcAAAQYBaYACwCGuQAE/+BAMQ8RNAoLGgs6BDgKSAVWC6oLvgvNC9kLCiELAQsDBwAfCy8LAi8LPwtPCwMLQBIWNAu6AqAAAwGstwICAQQHCAwIuAFYsy8HAQe4AmBADgJPAwEDGg0BABkM08IYK04Q9DwQ9nE8TfRd/QA/PD88EO39K11xPAEREjldMTABXSsTESEVBgICFyESEjdXA8F39oEB/vEH7cYEoQEFzHX+Sv4TwgEwAnj5AAMAU//mBBcFwAAYACQAMAENtTAIHR80Jrj/+EBsHR80xxHHE9cF1wcEdRB2FIQQAyYAKgw2ADsMRgBMDG4EYwhnEWgVdyeHJ5cNmBikDakYqRqmHqcnpiypMLkatx4XdxOGE4YUhycElwwBDJcAAQAcLpgMAQwrCZcAAQAlAy5AEhY0Py5PLgIuugKOABz/wEAQFhg0cByAHAKgHAEcHAYSKLj/wEAJEhY0MChAKAIouAKOQA0SDT8iTyICIkASFjQiuAKOQBoGBR/YCXcr2E8PAQ8aMhnYA3cl2BYZMdPCGCtOEPRN7fTtThD2cU3t9O0AP+0rXT/9XSsQETkvXXEr7V0rARESOV0REjldABESOV05XTEwAXFdAHFdKysBJiY1NDYzMhYVFAYHFhYVFAQjIicmNTQ2ExQWMzI2NTQmIyIGAxQWMzI2NTQmIyIGAUhtY+XT0edqYHp//v3XyIWddrlfT1BgX05RYBp3WVdydFlnZQMXLqFgpNbWpGafKjG8e8v+aXzYd8cBUVReX1RPX2D9PXSCfXZnfY4AAAIAQf/mBBQFwAAXACMA0EBYOxFLEWULegiJCKkFqQimDqYTtQC5A7UOuBG0E8UAyhHAExE0E1YLWQ1fEVITYBMGGQV3FpkX3RDfFAVoEwEABAEHGBIfGy8bAhtAEhY0G6YPBRAhICECIbj/wEAQEhY0IaYwCQFPCd8J8AkDCbgBT7OgAQEBuAEhtRAEIAQCBLj/wEAbEhY0BKYVDRjYTxIBEholAdgAdx7YDBkk08IYK04Q9E3t9O1OEPZxTe0AP/0rcfRd9l1x7StxP+0rcQEREjkAERI5MTABcV0AcV0TJRYWMzI2NwYjIgI1NAAzMgAREAAjIiYBNCYjIgYVFBYzMjZdARAKVEVXehFqn637AQnN3wEe/tbvrNQCXn1STmdwVFFvAVMeU1Cg/HsBC9bfARH+p/51/m7+nLcDHIiWe4yOhYAAAgAAAAAFvwW6AAcACgFBuQAH/9hACTc5NAYoNzk0B7j/wEAJKDU0BkAoNTQHuP/YQFAhJzQGKCEnNCkAKgQqBSgKLww4ADcFPwxqAGoCZQNmBWgIZwroAw9KBgECCAkBAwoJCQQHCQEBIAAHFAAABwYJBAQgBQYUBQUGCApAGh0+Crj/wEALGh00CiUCAwMGBAm4AbxADgYHAgUEBAEACAwXFxoAuAJhQAsfAQEgATABgAEDAbgCJEAJHwkBMAmACQIJugIkAAQCYUAJIAUBBRkLXmMYK04Q9F1N/Rn2XXH0XXEY/U5FZUTmAD88PBA8PzxN7RESOS88/SsrPIcFLiuHfcSHLhgrh33EBxA8PIfExLEGAkNUWLQJNAkNNAArWTEwAUuwC1NLsB5RWli5AAP//rIIBAq6//4AB//8sQYEODg4ODhZAXFdKysrKysrISEDIQMhASETAwMFv/6+gP22ef7GAjsBOSrKxgFN/rMFuvyKAiD94AAAAwCWAAAFYgW6ABMAIAAsANhAP3cqAWgOeCrmBPYEBAkhFQkGKCwhJRYSHxVPFQIwFa8VAhUVFCMiJRITCCAUJQEAAhsncAaABgIGSygnrwwBDLj/wLMJCzQMuAKMQCEwLkAuUC5gLnAugC6QLqAuCCAuMC4CLhQiIAAgEzATAhO4AouzLTFTGCtOEPRdPE39PE0QXXH2K3FN7fRd7QA/PP08Pzz9PBE5L11xQ1xYuQAV/4CyHTkVuP/Asho5Fbj/gLETOSsrK1k8/TwBERI5ABESOTEwAUuwC1NLsA9RWlixCiA4WQFdAF0TITIeAhUUBgcWFhUUBgYHBgUhAREzMjc2NjU0JicmIwMRITI3NjY1NCYmI5YCSq6rh1pvX4aQXaF2Sv7l/g0BKMKtKkxXS0os0aoBEqArQlNAecoFuh1cmV9nrCsnvH9kvXENCAIExv6tBQlXR0RVCQX9uf54CQxdTkJcKgAAAQBh/+cFXgXTABoA1kBOhgmJFIkWnwCYBscJ1APUC/UDCSUJKAwoDSkUKRZ1BXUJhgUIBxMHFxcTFxcpAioDJQUHKAWZBZcJyQPFCwU/AU8BAgFSEAAB4ADwAAIAuP/AsxEYNAC4/8CzCg00ALgBWkAXGC0ECA5ADhI0DktfDwFPDwEPQBUYNA+4AShAIhItCgMP7w5WAO8AAU8BAgEaMBwBHBUnoAcBDwcfBzAHAwe4AoyzG35TGCtOEPRdcU3tThBd9l1N7fTtAD/99CtdceQrP/30KytdceRdMTAAXQFdXV0BBQYEIyAAERAAISAXFhcFJiYjIgYREBYzMjYEPwEfQv7N7P7c/ogBegE0AQ2oZDL+2xqldqPLyKB2qgIbW/DpAY8BWgFuAZWfXrBGcoTq/vr+6uyWAAACAJQAAAVhBboAEAAfAH9AMygFKApHF2UEZQwFKhc5F0gWWRZoFgU5FzYbhxuZBZYLBR8RJQEAAhMSJQ8QCBknrwcBB7j/wLMJCzQHuAKMQBOAIQEgITAhAiEREiAAIBAwEAIQuAKLsyAxUxgrThD0XTxN/TxNEF1x9itxTe0APzz9PD88/TwxMABdcQFdEyEyFxYWEhUUBwYHBgcGIyEBETMyNz4CNTQmJicmI5QCHbdggbhgLTdmTYNipP3TASjdfDdIXzw8bFM+tQW6HCbC/ufOtYOgY0sqHwTC/DUOElbFqqq2ZhIOAAABAJUAAATwBboACwCQQD0IBQQHCCUGEh8FATAFrwUCBQUJAwQlAgECCgklCwAIBwZLAwJICgALAQsaIA0wDUANAw0ECSABIAAwAAIAuAKLswwxUxgrThD0XTxN/TxOEF32XTxN9Dz0PAA/PP08Pzz9PBE5L11xQ1xYuQAF/8CyHTkFuP+Asho5Bbj/gLETOSsrK1k8/TwDBRA8PDEwMxEhFSERIRUhESEVlQQ//OkC4P0gAzMFuvj+u/f+cfcAAQCXAAAEhAW6AAkAckA/CAUEBgUlByAIMAi/CN8IBC8IkAgCCAgAAwQlAgECCQAIBz8GTwYCBlIDAAIBAhogCzALAgsECSABIAAwAAIAuAKLswoxUxgrThD0XTxN/TxOEF32XTxN9F08AD88Pzz9PBI5L11xPP08AwUQPDwxMDMRIRUhESEVIRGXA+39OwJk/ZwFuvj+pfj9kQAAAQBi/+cFvQXTACAA2EBGOB5LHlYHdgh2DIUIhAyFF4QbCQYXBhsSFxIbKBEoGCgaKB4ISAtbBFQJWgtqBHsEehh0GrYOthDHDcYQ1xDnEA4DHAYgALj/wEAfGjkfAAEAJQIBARYcLQYJEkAOEjQSS08TARNAFRg0E7gBKEAqFi0PAwABASAZXxMBEycSVgIfICADAhogIjAiAiIZJ6AKAQ8KHwowCgMKuAKMsyF+nxgrThD0XXFN7U4QXfY8Tf08EPTtcRESOS88AD/99Ctd5Cs/7RE5Lzz9cSs8ERI5MTAAXQFdXQE1IREGBCMiJAI1NBI3NjMgBBcFJiYjIgYVEBIzMjY3NQM/An5d/p+15v6qrMC5jdIBEQEzLP7aH6uAwuXovF27QwIb9/24WonBAWfT5QFkX0nlyjdsffby/vv++0k0ugABAJYAAAUqBboACwCjQCUJBAUKAwIJCiUEEq8DAQMDAAYFBQIBAgcICAsACAUIIAbPBwEHuAKLQCJADVANYA0DcA2ADQIgDTANoA3ADQQNAgsgASAAMADAAAMAuAKLswwxdRgrThD0XTxN/TxNEF1xcvZdPE39PAA/PDwQPD88PBA8EjkvXUNcWLkAA//Ash05A7j/wLIaOQO4/8CxEzkrKytZPP08AwUQPDwQPDwxMDMRIREhESERIREhEZYBKAJEASj+2P28Bbr9vwJB+kYCgf1/AAEAjAAAAbQFugADAG+5AAX/wLMyNDQFuP/AsyMlNAW4/8BAPxQXNAAFQAVQBYAF4AUFHwVgBXAF8AUEgAUBAgECAwAIAgPZAQAAsADgAAPAAPAAAiAAMADQAOAABABuBDGfGCtOEPRdcXI8Tf08AD88PzwxMAFdcXIrKyszESERjAEoBbr6RgABAJkAAAXDBboACwGRQBoIBgESEgoKBQMCAwQGBgcJCgkICgUJCAkKCLgBt0ArBwYUBwcGAwQEIAUKFAUFCgoJAwMGCgMJAwgLBgYHBQQEAgECAAsLCAcIBLgCZLIFSAi4AmRAEgcaIA0wDQINAgsgASAAMAACALgCi7MMMWMYK04Q9F08Tf08GU4QXfYYTe307QA/PDwQPD88PBA8GRI5LwEREhc5ABIXOYcFLhgrBH0QxIcFLhgrCH0QxIcIEDwIxAMIEDwIPLEGAkNUWLUJIAsNNAO4/8qyCCc0ACsrWTEwAENYQBkmBicJkASYBqAEsATABAeEBqgE6AT2BQQJuP/gszdSNAm4/8BAJDdSNCUGPQp0A4YDmQOZCZoKqgO6A8kDCsED0AP8CgM9CkIDAnJxXSsBK3FdWUNcWLkABv/osxILPwa4/+hAEw8LPwQwDRY/BDAMFD8EIAsSPwO4/9CzDxk/A7j/0LMOFz8DuP/Qsw0WPwO4/9CzDBQ/A7j/0LMLEj8DuP/Qsg4TPwArKysrKysBKysrKytZAV0zESERASEBASEBBxGZASgCVgGO/dgCRv6B/m3wBbr9dQKL/cX8gQKw9f5FAAEAnQAABKUFrgAFAD1AGlAHAQIBAgQDJQUACAQFGgcCAyABIAAwAAIAuAKLswYxuRgrThD0XTxN/TxOEP48AD88Tf08PzwxMAFdMxEhESEVnQEoAuAFrvtJ9wAAAQCRAAAGGQW6AAwCGEALCwMmCCYLAwQDAQO4/4BACRw6NAogOjs0Cbj/4LM6OzQJuP/gQKQcLjQKIBwuNAYJCArjCewKBAQJCgoTAhwEEAkfCiMCLAQgCS8KZwJoBGUJagp3AngEpAmqCrUJugr2CfoKFp8EkAmfCsYJyQrXAtgE1gnZCucC6ATlCeoKDXcJeAqDAowEgwmMCpACB1gLZQJqBGcJaAp2AnkEB0QCSwRECUsKVwhXCVgKBxgKLw40AjoENAk7Cj8OBwMCDAQGCQkKFQIaBBcJB7EGAkNUWEAfAgQDCgkFDAcHMgYODDIAAAMQAwIIUAgNNAtQCA00A7j/gEAOCw00CEAOJzQLQA4nNAO4/5xAEA4nNAMLCAMBAAQBAgcKAAgAPzw8PzwREhc5KysrKysrXQEv7RDU7RESFzkbuP87QC0DCgkgBAgJCTIDBBQDAwQCCwoKMgMCFAMDAgsIAwMMBAICDAoKCQkHCB8OAQ64AQ2zBwYFBLoCOAAF/8CzW100Bbj/wEAXU1Q0BTIHQAd/CAEIvX8DAQO9CyALDAK4AjhAEgEAAEBbXTQAQFNUNAAyHwwBDLgBDbMNMXUYKxD0ce0rKxA87hA8GhkQ/XH9cTwaGBD9KyvuEDwQ5HEAPzwQPBA8PzwSFzmHBS4rh33Ehy4YK4d9xCtZMTABS7ATU1i5AAj/4LELIDg4WQFdXV1dXV1xcisrKysAK3FdMxEhAQEhESERASEBEZEBuwEKAQcBvP7t/t3+4/7eBbr8GAPo+kYEgvt+BIL7fgABAJgAAAUjBboACQHOQA4JAwYIGQMXCAQSCAIDA7j/ALMSCz8DuP/As1tdNAO4/8BAKlNUNAMyBwgUBwcIAwgCAgcDCQQCAgkHCAMEQFtdNARAU1Q0BDIGzwUBBbgCi0AZQAtQC2ALA3ALgAsCoAvACwIgCzALAgsICbj/wLNbXTQJuP/AQA5TUzQJMgEgADAAwAADALgCi7MKMXUYK04Q9F08Tf0rKzxNEF1dcXL2XTxN/SsrPAA/PD88ARESOTkAEjk5hy4rKysrh33EsQYCQ1RYuQAD/+BACQ4nNAggDic0A7j/wLcJDTQIQAkNNAArKysrWTEwQ1i5AAP/gLYLNQiACzUDuP/AQD0aLjQIUxouNAUDFgMyA0ADBEYDhQiQCKAIsgjkAwbEA88I2ggDIAMvCDQDOwhPCJIDnwigA68IsAO/CAsHuP/AQAkzNTQCQDM1NAe4/+BADS8yNAIgLzI0AgcUNQe4/5dACSEuNAJUIS40B7j/wEBGHiA0AlQeIDQIAgcHGAIDFwcsAicHOwIzB04CQAdcAlYHCRQCGwdNAkUHmgerB8sC2QLoAucH+QILJwIoB0oHeAeIB6wCBgFdcXJyKysrKysrKysrAF1dcXIrKysrWQBdMxEhAREhESEBEZgBIAJYARP+1/2xBbr8LQPT+kYDvPxEAAACAFn/5wXnBdMADwAbAKJAVZcFlwiYDJgOBAgBBw4IDwcYJxh4CXcSB3cReBWGBIkIiQyGDoUSiRSIFYgXiBiGGgwHEggUBxoVEhoUGhgVGgcTLQ0JGS0HAxYnrwoBAAoQCiAKAwq4AoxAIDAdQB1gHXAdgB2gHQYgHfAdAh0QJ6AAAQ8AHwAwAAMAuAKMsxx+wxgrThD0XXFN7U0QXXH2XXFN7QA/7T/tMTABXV1xAF0TNDc2Njc2MyAAERAAISAAARQSMzI2NTQmIyIGWUMyrWeJswFEAYX+fv69/rn+fgEx5rGx4923t+AC1OCYcLIrOv5u/pr+nf5vAY8BaPn+/////Pj7AAACAJUAAAT4BboADwAbAHdAJQYFuRS5GANHBQFnBdYFAhIRJQ0ODgAbECUCAQIPAAgWJ68HAQe4/8CzCQs0B7gCjEAWHx0wHWAdcB2AHQUdEA8gASAAMAACALgCi7McMVMYK04Q9F08Tf08TRBx9itxTe0APzw/PP08EjkvPP08MTAAXXEBXTMRISAXFhYVFAYGBwYjIxkCMzI2NjU0JicmI5UB2wEOUn6qYpdOasnBoq92Q15INaAFuhYh3a+HuGkRFf3XBML+YC5iQVBoDQoAAgCWAAAFvAW6ABUAIQD4QII5D0kPVwdqC2oMqgmnDqAjtg7YCQoGCAYKFwgWCjYORg5GDwcIEAkRFA4UDxQQNg42D0cPdQ55ENMKC3gJeBl2HYgJiBmGHQYJFhQJDA8OUw51DoQOlA6jDgUOIA0MFA0NDA8MFQ0XFiUTEBQBYBSgFAIUFAAgISUCAQINDg4VAAgOuAG8QCcADRANAg3UGyegBrAGwAbQBgQGh3AjASAjMCMCIyEVIAEgADAAAgC4AouzIjFjGCtOEPRdPE39PBBdcfZd7fRd7QA/PDwQPD88/TwSOS9dcTz9PAEREjk5hy4rXQ59EMQBETkAERI5MTAAXQFxXV0zESEyFhYVFAYHFhYXEyEDLgIjIxERMzI2NjU0JicmIyOWAm/r1YDCwWB9arP+ntZyVF5mPNvVajxPSCS05wW6T8qCpdccOIar/uIBP6tZIf2cA04kWEJKWwwFAAABAEr/5gTyBdMALAHQQD25EbgdtijGLAQHEwcVFxMXFRgrZQVlKHQGeA10KNkM1iMMWQpVDlUiWSNoDGYSZyFpKGcsdx2GHZYhDBIjuP/gsx4fNCO4/+BAZRkaNFEiUSPBIsEjBHEicSOBIoEj4SLhIwYrCioNJCIkIzkNNCNLCksNRCJDI2oNZSN5DXoiiQ2KIqYKpw2oIhMJCgkNBiIGIxkKGQ0WIgciIwoNBAEXVhhAGSA0bxgBbxifGAIYugJlABv/wEAMGjkfGwEbLRQDAEgBuP/AQEkaIDQwAUABUAFgAZABoAGwAcABCAHuBEAaORAEAQQtKgkY7/8XARdAExc0F0sHJyYaLh8noBCwEAIQSwHvESAAMAACABkt0lMYK04Q9F1LU1ixAEA4WU3t9F3tThD2Te30K3LtAD/9cSv0XSvkP/1xK/RdcivkEhc5XV1xcisrQ1xYuQAi/+CzGx0+I7j/0LMbHT4juP/jshM5Irj/4LITOSO4/8myEjkiuP/QQA8SOQ0gEjkKIBI5CiAPOSK4/+hADgw5DSANOQoYDTkKGBM5KysrKysrKysrKysrK1mxBgJDVFhAFToKOg01IjUjSwpJDUMiRiOmCqkiCgBdWTEwAF1xAV0TJRYWMzI2NTQmJyYnJicmNTQ2NjMgBBcFJiYjIgcGFRQXFgQWFhUUBgQjIABKASAan4ePkT1MNLnuYId/76kBFAEXB/7YE319gUkvLDgBsM91jP8Av/7q/tYB3RyRiHlRNEkbEi47VnmucMNm8soNcWM1Ijk0JS9mbb2LftxrAQEAAAEALAAABLkFugAHAHJAIy8JMAQwBVAJcAmACZAJBwYBBQIlBAMCBwAICRcXGgR/BQEFuAEtQAoGByABMAB/AAIAuAEtQBEDDlACcAKAApACBAIZCP2sGCtOEPRdS1FYsQJAOFk8TfRdPP089F08RWVE5AA/PD88/Tw8PDEwAV0hESE1IRUhEQHf/k0Ejf5OBML4+Ps+AAEAk//nBSQFugAZAIpAOAcIBwkHEBcIFglHCEcJB1cJVhCWEJcRmBWbFqcQtxbXFeUG9gYLDQwMAQACByUTCQwLIA3PDgEOuAKLQCJAG1AbYBsDcBuAGwIgGzAboBvAGwQbAQIgACAZMBnAGQMZuAKLsxoxdRgrThD0XTxN/TxNEF1xcvZdPE39PAA/7T88PBA8MTABXXETIREUFxYWMzI2NjURIREQDgIjIiYmJyY1kwEoCxOPfH6AGgEoMIHYrtLZfhQdBbr85r04Wm1nlq4DK/z+/vjalllhm1V+9gAAAf/9AAAFWAW6AAgAxbkABP++QD4LNcAKAQQDBAUDBwQFBAMFAQQDBAUDIAIBFAICAQQFBAMFIAYHFAYGBwEEBwMGCAcEAQMCAwkEAAUKCAFWB7gCZ0ALBgYFBQMDAgIACAq7AhcACAAGAhe1BwcIIAACuAIXtwEBIAAwAAIAuAJmswleYxgrEPZdPBkQ5BgQ/TwZEOQYEOQAPz88EDwQPBD25AEREjkSORE5ABEXORESFzmHBS4rCH0QxIcFLhgrCH0QxAcIEDyHCBDEMTABXQArIREBIQEBIQERAhb95wFbAVkBUgFV/eUCaQNR/bwCRPyt/ZkAAQCS/mMChAW6AAcAUEAyBjAFQAUCBTcAAz8ETwQCBDcBEAASAwIGAgcEBRAHAQf0BZsAACABMAHQAQMBYAhnfBgrEPZdPBDt7V0QPBA8PBA8AD8//V08EP1dPDEwExEhFSMRMxWSAfLn5/5jB1fd+mPdAAACAEn/6AQuBD4AIwAyAXFAaAcaCBwFHRYaShtIHEkl2xDfEQk2GUYZVyZmGWcmhiaSGZMaphq5G8cayBsMBgYNFRYGGRYnBikVWRl3AoYCpga1BsYGDL802RACHSQyMREsDSRAKy40JEAiKDQkQBkdNG8k/CQCJEYduP/AQDAODzQ9HQEAHRAdsB35HQQdHSwBMwBADg80DwAfAAIAVSFAHBE/IUAbED8hQBgaNCG4AnS1BAcMDQosuP/AsxwRPyy4/8CzGxA/LLj/wLMYGjQsuAJ0QEAUCx4xJggpCSgNWR8MnwwCHwwB/wwBDEAOFjQMGk80ATRgAAEAjjABAQEzKSFfFwHfFwFPF18XbxcDFxkzaUEYK04Q9F1xck3t9HHtXU4QXfYrXXFyTe305P08AD/tKysrPzw//SsrK/RdK+QSOS9dcSuxBgJDVFiyLx0BcVntsQYCQ1RYuQAk/8C3Gx00VCRkJAJdK1ldKysrERI5Aw4QPDw8MTABcV0AXXEBJzY2MzIWFhUDFBYXISYnJicGBiMiJjU0NjY3Njc1NCYjIgYBBgYHBhUUFjMyNzY3NjUBZf8r0s+8uEsDGyX+6gsQBwNIpF2kvVabksVMUG9LVAFeNuokN1hETEUzEAsC4i6alFmJt/64jIVMHDcZCEZGsohajUscJSAcUUU7/tISMhgnPDtWMiY3JGUAAgCH/+gElAW6AA8AHACduQAS//hAMQs5NxtHGwISVgZWClYWVhhZHPcHBjUEOw07EzUbRQRLDUsTRRuUB5kJCgwOAQIBABq4AnSyBQcUuAJ0QBMLCw8AChchCBpwHgEeECkCAyYPuAEpQAwBcACAAAIAGR0/QRgrThD0cTxN7f085k4QcfZN7QA/PD/tP+0/PDEwAHFdAV1DWEALZgZmCmYWZhhpHAVdWQBdKzMRIRE2MzISERAAIyImJxUTFBcWMzI2NTQmIyIGhwEZgrLC/v79uVuxQBI0SXldg4RnZYYFuv3wlP7n/vn+8P7aW1mcAiqlT3Cfq7ahnQAAAQBV/+gEPwQ+ABkA4UBRWA9ZElkWaA9pEmkWfRh5GZcClwzGEMYY1xDWGOkG6QjpE+kV+AYTOBM4FUoSShZGGFkMaQwHOhI3FjcYA3cFdw+HBYYPiRmoEqcWuRK2FgkOuP/AsxgbNA64/8C1EhQ0DjMNuP/AsxkeNA24/8CzDxE0DboBBAAKAnRAEhELAEAYGzQAQBIUNAAzkAEBAboBAQAEAnRAIBcHAUASFDQBIQAvDUASFDQNIU8OAQ4aGwchFBkaWEEYK04Q9E3tThD2XU3tK/TtKwA//fRd5CsrP/30KyvkKysxMABdcQFxXQEFJiYjIgYVFBYzMjY3BQYGIyIAERAAMzIWBDH+6w5jT2l9f2tQZhUBFCv0zen+6wEW7cLlAuwyU1SRqr2cW28vvsIBJgEEAQcBJacAAAIAVP/oBGEFugAPABwAkEAtElkGWQpZElYWVhhZHJgHmQn4CQlwHoAeAjoDNAw6FTQZSgNEDEoVRBmZCQkUuAJ0sgULGrgCdEAOCwcODwABAAoXKQ4NJgG4ASlADw8AGo8eAR4QIQgZHVg8GCtOEPRN7U4QcfY8Te39POYAPzw/PD/tP+0xMABdAXFdQ1hADWkGaQppEmYWZhhpHAZdWSEhNQYGIyIAERASMzIXESEBFBcWMzI2NTQmIyIGBGH++0GxWrf++/7CsoIBGf0SL0R6YYiEZ2SHnFtZAScBCAEOARmUAhD8cKpMbqWkt6GfAAIAQf/oBCcEPgAUABwBo7kAEP/4QEYLOZkJmg2WEKgFpwq7CbsNuBoICBQBSAJHBkYKTx6oDbYGthrHCsgM1grYDPgH9w0NHA8cFUAbHTQVQA4RNA8VvxXPFQMVuP/Asw8ePxW4/8CzDhc/FbgCjUAMDw4SUA5gDgIOGBIBuP/AthkbNAEzEgC4/8CzHSA0ALj/wLMiKTQAuP/AsystNAC4/8CzGBw0ALj/wEAPDg80oAABAAAQAAIAXxISuAJ0swQLEhi4AnRAJAsHACEBLxUhTw4BDhovHl8ebx6fHgQeDyEIQA0PNAgZHWlBGCtOEPQrTe1OEF32XU3t9O0AP+1DXFhAFBhAKBQ/GEAeDz8YQBsQPxhAHBE/KysrK1k//UNcWLkAEv/AsygUPxK4/8CzHg8/Erj/wLMbED8SuP/AshwRPysrKytZ9F1xKysrKytDXFi5AAD/wLISOQC4/8CyFzkAuP+wswkKPgC4/8CyQSE/KwArKytZ5CsREjldQ1xYQBQOQA8ePw5AHBE/DkAbED8OQA4XPwArKysrWS88/SsrcisrPAERMzEwAV1xAF0rAQUGBiMgJyY1EAAzMgADIRYWMzI2EyYmIyIHBhcC+gEYNumv/uuFaQEU0+0BEgb9QAOCYUJaJwN4Vlw8PAEBUi+aobWR3QEIASv+x/69fYtIAWx6f0NDcwAAAQAYAAAC5gXTABYAuEAyNgQBKgQgECARWQSAGAUIBL8YAhUWEQIUEhYRDhMPABAOEwEAEAIUCQgPCwFfC/8LAgu4AnRACgYBEQ8WAf8WARa4AnRAHhAAAAHwAAEABhMUCgkzPwhPCFAIAwgoEC8RXxECEbgBBEANDhMmAhRfAKAWwBYCFrj/wLYJDDQWGRd4uQJpABgrThD0K3E8Tfw8/Tz8XTz0XRnkABg/PD9dcTz9XXE8P/1dcTkyDw8PDzEwAXFdAF0TMzU0NjYzMhcHJiMiBhUVMxUjESERIxicOZl1eHMmQz49NdLS/uecBCZQhoRTJMQQOVFL3fy3A0kAAAIAVP5RBGAEPgAjAC8BTkBidx2HHQISDA1wMYYNgDEEIAEjAiMDMAEzAjMDQAFDAkMDWw9ZFFklVilWK1kvaw/4EfgTEjsNMxY7KDMsSw1EFksoRCzwDP0XCo4MAQwLDA0LKgwNJw4WFxUtDQwXFgQYJAG4/8C1GRs0ATMAuP/Asw4RPgC4/8CzCww+ALj/wLMoKjQAuP/AsyMlNAC4/8CzMTQ0ALj/wEAJFRs0YAABAF8FuAJ0sh8PJ7gCdLIOCi24AnRACxUHGBkGKikLJhoYuAEpQAkZGRoajzEBMQG4AbhACgAzJCESGTBYPBgrThD0Te307U4QcfY8TRDtEP3kAD88P+0/7T/99HIrKysrKyuxBgJDVFi5AAD/wLMOETQAuP/AsgkMNCsrWeQrARESFzkAERI5ORESOTkHCBA8MTAAcV0BXXFDWEANaQ9pFGklZylmK2kvBl1ZAF0XBRYXFjMyNzY3NjU1BiMiJyY1EAAzMhc1IREUDgIjICY1NBMUFjMyNjU0JiMiBnkBQQgdKFZuNyUTDX7A1n1iAQG/xYABBz5wu4/+8uL8g2BnjohoZYNGJzgVHiEWMSNem6y1j9UBCwEarZX8R7y6ajy5jg4Cg6mdoZ6loJ0AAQCSAAAEWQW6ABYAskArDwEfATkBMwIzEEIBQhHeAfkBCQcFFgUkAlgRaBEFAQECExQREhMDFAIBD7gCdEAdAwcJCgoUFQoWAAALCiYICUAgJDSvCQH/CQEJGhi4/8BAFiIkNJAYoBgCcBjwGALvGAEYABQmFhW4/8BADyAkNKAVAfAVARUZFz88GCtOEPRxcis8Tf08ThBdcXIr9nFyKzxN/TwAPzw/PDwQPD/tOTkRFzkDDhA8CDwxMAFdAF0BETYzMh4CFREhETQmJiMiBgYVESERAauIvWGcTx3+5yBRPUZuM/7nBbr95Z9IcIiP/ZECMadaNUSJhv3sBboAAAIAkwAAAawFugADAAcAd7kACf/AQD8RCj9ACVAJAoAJsAnACdAJ7wkFHwlgCX8JoAmwCQUDBgcABQQDDwABQADQAOAAAwBdAgEABgUGBwQKAgcmAQS4/8BACSEkNAQZCD88GCtOEPQrPE39PAA/PD88Pzz9XXE8AwUQPDwQPDwxMAFxXXIrExEhEQERIRGTARn+5wEZBLYBBP78+0oEJvvaAAEAkwAAAawFugADAFO5AAX/wEApEQo/QAVQBQKABbAFwAXQBe8FBR8FYAV/BaAFsAUFAgEAAwAKAgMmAQC4/8BACSEkNAAZBD88GCtOEPQrPE39PAA/PD88MTABcV1yKzMRIRGTARkFuvpGAAEAfgAABpgEPgAnATu5ACn/wEBdEQo/BQYGDBUGFgw0AzQINBg0I0QCRQhFGEQjDCADLylTCWApgCmfKaQGpwemDLUGtQywKdAp4CkOACkvKVApnym/Kd8pBilAGhw0PylQKYAp0CngKQUHIQQHGh0WuAJ0sgoHIbgCdEAeBAcQEREnGxwcJicKAQAGDxAmEhFAWjVgEQFvEQERuAJGQA8aGyYdHEBaNW8cAWAcARy4Aka0JSYmJwG4ASmyAAAnuP/Asw8JPye4/8BANhEKPydAWjUnQEE1J0A8NSdAJCc0J0A6PTQvJ88n3ycDDycfJ4AnAwAnICcwJ/8nBCcZKOM8GCtOEPRdcXIrKysrKysrPE0Q7RD9PPZdcSs8/Tz2cV0rPP08AD88Pzw8EDwQPBA8P+0/7QEREjkAERI5MTABcitxXQBdASsTIRU2MzIWFzY2MzIWFxYVESERNCcmIyIGBhURIRE0JiYjIgYGFREhfgEDi8BmljBGolx1oigd/ucdJ1E7aC7+5x4/NkFoLf7nBCaRqVRVVVRfXESY/VkCX54uPEiLlv4CAkabWixGhJn9/AABAJEAAARZBD4AFgCfQBgHExcTWghoCAS4BAE0CDQQRAhED+kQBQa4AnRAHREHDg0GDAsLAQAKAgEmFgBAICQ0rwAB/wABABoYuP/AQBYiJDSQGKAYAnAY8BgC7xgBGAoLJgwOuAEpsg0NDLj/wEAPICQ0oAwB8AwBDBkXPzwYK04Q9HFyKzxNEO0Q/TxOEF1xciv2cXIrPE39PAA/PDwQPD88P+0xMABdAXFdISERNCYmIyIGBhURIREhFTYzMh4CFQRZ/uckUTlJdCv+5wEFi9Ndmk8fAh6sZThQhLL+HwQmnLRDaIR7AAACAFL/6ASaBD4ADQAZAJdASOgB5wj3E/cVBMcC6AUCEhkFGQkCWRBWE1YWWRiXApgGmAiXDLgJ1QLbBdwJ1QznBecG6A0QpwjLAswGwwjGDAV1CIkGhAgDEbgCdLIKCxe4AnRAFAQHFDkHGmAbcBsCGw4hABkaWEEYK04Q9E3tThBx9k3tAD/tP+0xMABxXQFdcUNYQAlpEGYSZhZpGAQBXVkAXQFdEzQSNjMyABUUACMiJCYlFBYzMjY1NCYjIgZSiv2c8QE0/snskv73igEglm5ulZVubpYCIowBBor+x+/x/sOE/6ieqKignKioAAACAIv+bASXBD4AEAAcAJpALjgTSBMCEjQDOQ05EzQbRANJDUkTRBv5GwlWBlYKWRJWFlYYWRz2B/kbCAEABhq4AnSyBQcUuAJ0QBYLCxAPDhchCBpwHgEeESkODg8mEBABuAEpQAtwAIAAAgAZHT9BGCtOEPRxTe08EP08EOROEHH2Te0APzw/7T/tPzwxMAFdAF0BQ1hADWYGZgppEmYWZhhpHAZdWQBdEyEVNjYzMgAREAAjIiYnESEBFBYzMjY1NCYjIgaLAQYzrmq5AQL+/LlYj0/+5wEWjmZigoZjZ4gEJpxQZP7e/v3+9v7ZRlX96QO5s6uds6einwABAIcAAAM3BD4AEACoQCiXBQEJDgFTBWYFdQUDLxJYDmgOcBIECgkPDB8MAo8M/wwCPwxPDAIMuAJ3QCkHBwEACgMCBgooAAkQCTAJcAkECRp/Ep8SAl8SfxKvEtASBBIQACYBA7gBKUALAgKAAaABAgEZET+5ARwAGCtOEPRxPE0Q7RD9PE4QXXH2XRlN5AAYPzw/PD/tXXFyOTIxMAFdAF1xAEuwF1NLsDVRWlixCjI4WQBdISERIRU2NjMyFwcmIyIGBhEBoP7nAQVDa0RgWVdHPTtSLwQml2tENfUuQar+8QABADD/6AQQBD4AKgLCQMAGEQYjCCcXERcjmBKYFJcnlSoJBxRGFAISuw25Dsch5SP4DfYiBikNVQ1lDZULlxKnIrkMB0EjQCREJmciZCaHEocUhiKDJAk3JkUGRgtKDU8PRiFCIgciJCcmNww1ITUiNSM1JAcGCgURCSEYDScMIiIiIwckIkAscwx4FHkVdil1KogVhCqaFZUqtCK0Iw2AAY8XjBiZKqkqsCwGFyEWQCEjNBZAHB80HxYB3xYBFjMIIVAljyUCJUAYHTQlGiy4/8BAFxEKP1AsATAsAS8sASweITAQARAzASEAuP/Asw8JPwC4/8CzEQo/ALj/wEAJCQ00ABkreLgYK04Q/CsrK03t9HHtThBdcXIr9itxTe30cXIrK+0AsQYCQ1RYQDUGAQEGARYBJiI2IUYhVAFZF2QBaRf2AQoBFwIEGiEiAigTDQwCKBpfBAEERigLUBoBGkYTBz/9XT/9XRESFzkREhc5ERIXOV1xG7kAIv/LsygqNCG4/8uzKCo0Irj/4LMeJDQhuP/gsx8kNCK4/+CzGRo0Ibj/4EAbGRo0aw0BNiJGIpgNlCLEItQiBiEiDA0EBBoAuP/AtRkbNAAzAbj/wLMXLT8BuP+wswkKPgG4/8CzIiU0Abj/wEAdGhw0AAEwAUABUAEEYAGAAfABAwABEAFQAWABBAG4/8CzExY0AbgBAUBNAAQBXwTwBAIERigLFkAZGzQWMxdAFy0/F0AJCj4XQDU3NBdAKy40F0AlKTQXQBocNA8XHxdfF28XBBdVGkAiJDQPGgFQGv8aAhpGEwc//V1xK/RdKysrKysr5Cs//V1x9CtdcXIrKysr5CsREhc5XXErKysrKytZMTABcV0AcXFxcV1dQ1xYuQAk/8lACQsSPw8oCxI/Ibj/7LYNOQwUDDkhuP/ssgw5Irj/6rELOQArKysrASsrWQBxXRMlFhYzMjc2NTQnJickJyY1NDYzMhYXBSYmIyIHBhUUFxYEFxYVFAYjIiYwARoSbmNtNyUUFUn+rFt+2uXa1Cj+9xFfWG8wIBwmAcFZWPTv2f0BLytSVSgcLyAVFBFLPlaZiryOizE+Qh8WIx4VHGZKS4aS0rAAAQAf/+gCkQWdABkAzUApIAAgASMKKQ86DkoOWQ8HGRUAGAMWFQAXEhMUARcSAhQBGAMJBwoHDBi4AQFADwAXoBewFwNgF6AXwBcDF7gBBLIVARS4AnSzABUGB7gCdEAODAsJLwovAAAvAV8BAgG4AQRAKBgDJhcSVRU/FJ8UrxQDYBSAFJAU0BTwFAUAFBAUIBQwFAQUGRp4oBgrThD0XXFyS7A3U0uwO1FaWLkAFP/AOFk8Tfw8/Tz0XTwQ9BnkABg/7T88/TwQ9F1x5BESOREzDw8PDzEwAV0BFSMRFBYWMzI3FwYjIiYmJyY1ESM1MzUlEQJ6wAsnHCdKGGJ8THo5CwmBgQEaBCbg/lSCKxwb2iozUUUxlQHP4NOk/okAAQCN/+gEUwQmABYAnEAXVxFnEZYFAwkGGQY8AjwRSwJLEecCBw+4AnRAEQQLFgAKFRQUCgkGExQmFRUAuAEpQA4WQCAkNK8WAf8WARYaGLj/wEAWIiQ0kBigGAJwGPAYAu8YARgKCyYJCLj/wEAPICQ0oAgB8AgBCBkXPzwYK04Q9HFyKzxN/TxOEF1xciv2cXIrTe08EP08AD88PBA8Pzw/7TEwAF0BXSE1BgYjIiYmNREhERQWFjMyNjY1ESERA046vWlrqkwBGR9SP0hyKgEZn1ViXqqWAqD+GOBlO0915AHA+9oAAAEACwAABFoEJgALARtAFQUoGi80BygaLzQGKBovNAgoGi80A7j/2LMaLzQEuP/AQCAaOjSaBAEGAwsICAoMCxUBFQISAxoJGgoiAC0LxwsMALj/8EAWHSA0CgAFCxQAGQslACoLNAA6C4cACbEGAkNUWLQKAQ0MBLj/wEALCRc0BAEACQEGAAoAPz88ERI5KwEREjk5G0ASCwAKBAsKCQkCAgEGCwAKCTkNuP/AQBgcKDQLDR8NMA1ADQQNFxcaEAo/Ck8KAwq4AjBACwQCOQsEPwRPBAMEugIwAAH/gEAPDDUAASABQAEDARkMxKAYKxlOEPRdKxhN7V3tEP1dGU5FZUTmXSsYTe0APzw/PBA8EDwSOQESOTlZMTABcStdAF0rASsrKysrIQEhExc2NzY3EyEBAbf+VAEnyDoXBg4QygEh/loEJv3itUUWLS0CHvvaAAABAAkAAAY4BCYADAHdQDEACwEKAAYCCgcFCRsAFgIeBBEFGgcUCR4KEQwMEisDKwYjCzkDOQZIA0gGmAOYBgkOuP/AQHcsRzQKAAsEBAUECQsKBAwbABoEFgUUCRkKFQwMIwAoBCcFLQkoCicMMQA3BT4JRgBHAkcFSAdJCXcAeAR3BXgJeAp3DIcAiASHBYgJiAqHDNkA2QTVBdUJ2QrVDOoA6gTkBeQJ6grkDPkA+QT2BfgH9gn5CvYMLbEGAkNUWLQIAQ4NBrj/wLMJITQDuP/AQBUJITQLQAkhNAMLBgMAAQcEAQYJAAoAPzw/PDwREhc5KysrARESOTkbtMILBAUguP9NswYKCSC4/0xAMgMADCALBgMDDAACAQQMAwUKCwcJCAYIBwcFBQQEAgIBBgwKCgkJAAovDj8OAg4XFxoIQQkBDgAgAAYCbQALAm0AQAADAQ60IAEZDcS5ARoAGCtOEPQaGU39Ghj9/RoZ/RhORWVE5l0APzwQPBA8PzwQPBA8EDwQPAEREjk5Ejk5ETk5Ejk5ABEXOSsrK1kxMAFdcSsAXUNcWLQLQA05Brj/+LINOQO4//i2DTkLQAw5Brj/8LIMOQO4//CyDDkGuP/gsgs5A7j/4LELOQArKysrKysrK1kBXQBdIQEhExMhExMhASEDAwFZ/rABEce3AQ+xywEV/qv+8re0BCb9SAK4/UgCuPvaAqv9VQABAAwAAARgBCYACwGYQIsoB8gEApgHuQHcAdUH8A0FCAcaBBgGKAY3ADgISAFZAXwBdQcKJgErBzYBOgdGAUoHmAv4BvgHCSUEJgcqCjQEOgpDBE4KwwQITApUBFkKZARtCngBfQqUBJYHugrVBNwK/AoNAwQHBwkKFgQgBCoKMwQ/CkYECRUEGQo6Ck4KawqnBLcEyQr2BAkHuP/wsxIYNAS4/9izFRc0BLj/4EAVDBE0AQQKBwQAAgEECgcECAAJCAMDuP/gtiktNP8DAQO4/+BADxYkNAMmAgkUAgIJBQYLC7j/4LYpLTTwCwELuP/gQBcWJDQLJgAFFAAABQYFBQMCBggJCQsABbgCbbIGMwm4Am1ACwhlTw2fDeANAw0DuAJtsgIzC7gCbUAS8AABAAAQACAAMAAEAGUMxKAYKxlOEPRdcRhN7fTtGU0QXfYYTe307QAvPDwQPD88PBA8hwUuKytxK4d9xIcuGCsrcSuHfcQBERIXOQAREhc5sQYCQ1RYtQogCSE0BLj/4LIJITQAKytZMTAAKysrXXFxcgFdcXFyMwEBIRMTIQEBIQMDDAF//pEBV7zGAUr+mAGJ/qfY2gIjAgP+3AEk/gn90QFJ/rcAAAEADv5RBFIEJgATATS0EigFARO4/+BAGAwPNAgWDQ80BxYNDzQGFg0PNAUWDA80Arj/wEAfGjo0BQYGBA0LDgYQAgATBgQTAgQDAwEBAAYTYBABELgBr0ASCw8NLw4oACAVMBVgFQPwFQEVuP/AsyImNBW4/8BAEhweNBUXFxoEOQNAGBk0fwMBA7gBJ0AJAkAYGTR/AgECuAEnQBIBOQBAHDY0IAAwAAIAGRTEoBgrThD0XStN/Rn0XSv0XSsY/U5FZUTmKytxck0Q9OQAP+1dLz88EDwQPAESORE5ABESORI5ORE5Bw4QPDEwACsBKysrKytdS7AQU0uwOlFaWLIEEAC6//AAAf/wsQMQATg4ODhZQ1xYuQAF/+hADg0RPxMQExk/ExASGD8FuP/wsxMZPwW4//CyEhg/ASsrKysrWRMhExMhAQcOAyMiJycWMzI2Nw4BK/74ASP+iUMlQ1d/UFFOGUI1Yl4ZBCb9DgLy/AK5XWI9IhHcDXNZAAAAAAEAAAAFOFIAAAAAXw889Qg5CAAAAAAAouM8HQAAAADSlH8b+vr8/RAACCQAAAAJAAEAAQAAAAAAAQAABz7+TgBDEAD6+vp6EAAAAQAAAAAAAAAAAAAAAAAADV0GAAEAAAAAAAI5AAACOQAAAqoAuAPLAHAEcwASBHMARgcdAFkFxwBaAecAXAKqAGsCqgBDAx0AHASsAFUCOQB1AqoAcwI5AJMCOf/9BHMAVgRzAKIEcwAzBHMATQRzACYEcwBbBHMAVwRzAFcEcwBTBHMAQQKqAMkCqgCqBKwAXwSsAFUErABfBOMAagfNAD0FxwAABccAlgXHAGEFxwCUBVYAlQTjAJcGOQBiBccAlgI5AIwEcwAjBccAmQTjAJ0GqgCRBccAmAY5AFkFVgCVBjkAWQXHAJYFVgBKBOMALAXHAJMFVv//B40ABwVWAAAFVv/9BOMAFgKqAJICOf/9AqoAJgSsAHMEc//tAqoAKgRzAEkE4wCHBHMAVQTjAFQEcwBBAqoAGATjAFQE4wCSAjkAkwI5/6IEcwCJAjkAkwcdAH4E4wCRBOMAUgTjAIsE4wBbAx0AhwRzADACqgAfBOMAjQRzAAsGOQAJBHMADARzAA4EAAAiAx0APAI9ALADHQAtBKwAQwXHAAAFxwAABccAYQVWAJUFxwCYBjkAWQXHAJMEcwBJBHMASQRzAEkEcwBJBHMASQRzAEkEcwBVBHMAQQRzAEEEcwBBBHMAQQI5AJICOf/pAjn/zQI5/9AE4wCRBOMAUgTjAFIE4wBSBOMAUgTjAFIE4wCNBOMAjQTjAI0E4wCNBHMARAMzAFYEcwBUBHMADQRzADsCzQBCBHP//gTjAIsF5f/3BeX/9wgAANgCqgC7AqoABQRkADEIAP+qBjkAPwW0AJgEZAAyBGQAPARkADwEcwABBJwAbwP0ACwFtAB6BpYAoQRkAAACMQAAAvYAJQLsABoGJQA3Bx0AWATjAFcE4wBlAqoAwwSsAFUEZABUBHP/7ARkAB8E5QAaBHMAYARzAGoIAADJBccAAAXHAAAGOQBZCAAASAeNAFgEc//8CAAAAAQAAIQEAABpAjkAmAI5AHIEZAAxA/QALwRzAA4FVv/3AVb+qQRz/+ACqgBLAqoASwTjAB8E4wAfBHMARAI5AJMCOQB1BAAAcQgAAAEFxwAABVYAlQXHAAAFVgCVBVYAlQI5AGoCOf+uAjn/vwI5/8EGOQBZBjkAWQY5AFkFxwCTBccAkwXHAJMCOQCTAqoAAwKq//MCqgATAqoAGgKqAM0CqgCRAqoAJgKqAGACqgA5AqoAAwTjAAoCOQAKBVYASgRzADAE4wAWBAAAIgI9ALAFx//9BOMAUwVW//cEcwAOBVYAlQTjAIsErABVBKwAbQKqAFsCqgAZAqoAKAasAFwGrABcBqwAKARzAAAGOQBiBOMAVAI5AIwFVgBKBHMAMAXHAGEEcwBVBccAYQRzAFUE4wBUBGv/7QKqAMgFxwAABHMASQXHAAAEcwBJBccAlAXAAFEFx//9BVYAlQRzAEEFVgCVBHMAQQTjAJ0COQB5BOMAnQMVAJUE4wCaA9UAkwXHAJgE4wCRBccAmATjAJEGOQBZBOMAUgXHAJYDHQCHBccAlgMdAFAFVgBKBHMAMATjACwCqgAfBOMALAPVAB4FxwCTBOMAjQXHAJME4wCNBOMAFgQAACIE4wAWBAAAIgTPAJoGOQBWBpEAVgTrAE4E2gBOA8wATgV5AE4DkgAwBbkATgRr/+0E1QC4AysATwjAACkIAABPBAAAmQgAAE8EAACZCAAATwQAAJgEAACYB9UBagXHAI8EqwBVBNUAnQSsAFUE1QIiBNUBBQWr/+kFAAHJBasCfgWr/+kFqwJ+Bav/6QWrAn4Fq//pBav/6QWr/+kFq//pBav/6QWrAcAFqwJ+BasBwAWrAcAFq//pBav/6QWr/+kFqwJ+BasBwAWrAcAFq//pBav/6QWr/+kFqwJ+BasBwAWrAcAFq//pBav/6QWr/+kFq//pBav/6QWr/+kFq//pBav/6QWr/+kFq//pBav/6QWr/+kFq//pBav/6QWr/+kFq//pBasC1gWrAGYFq//qBdX//wTVAJIIAAAAB+sBMAfrASAH6wEwB+sBIATVALIE1QCABNUAKggrAZgIawG4B1UAEAYAAPQGAABvBEAAOgVAADcEwAA/BBUAQAQAACUGAABVBkcAjARzAJAFq//HAesAjQPVAIYHFQAjA+kAGATVAJIC1gBcAtYAXATVALIC1gBNBccAAARzAEkFxwBhBHMAVQXHAGEEcwBVBVYAlQRzAEEFVgCVBHMAQQVWAJUEcwBBBjkAYgTjAFQGOQBiBOMAVAY5AGIE4wBUBccAlgTjAJIFxwAFBOMAGQI5/7oCOf+7Ajn/2gI5/9oCOf/hAjn/4gI5AEgCOQBHBHMAIwI5/6IFxwCZBHMAiQRzAI0E4wCdAjn/7QXHAJgE4wCRBckAnATjAI4GOQBZBOMAUgY5AFkE4wBSBccAlgMdACoFVgBKBHMAMATjACwCqgAHBccAkwTjAI0FxwCTBOMAjQXHAJME4wCNBccAkwTjAI0HjQAHBjkACQVW//0EcwAOAjkAjQXHAAAEcwBJCAD/qgcdAFgGOQA/BOMAVwKqAMkHjQAHBjkACQeNAAcGOQAJB40ABwY5AAkFVv/9BHMADgI5AJUCqv/XBHMADQTNAFoGrABcBqwAKQasADAGrAAvAqoAvAKqACYCqgC7A7j/9AXH/+gG0/+7Bz//uwPK/7sGmf+mB2v/yAa0/5wCOf8pBccAAAXHAJYFwAAABVYAlQTjABYFxwCWAjkAjAXHAJkFVgAABqoAkQXHAJgFJgBmBjkAWQXHAJoFVgCVBM0AWgTjACwFVv/9BVYAAAZ5AFYGagBiAjn/zAVW//8E6wBOA5wATgTjAI4COQCCBKgAbATiAJAEcwAPA68ATgTjAI4EUwBOAjkAkwR2AI4EcwAPBOUAkARzAAsDkABOBOMAUgTzAHYEKQBOBKgAdgSbABEGBwB2BsIATgI5/80EqAB2BOMATgSoAHYGwgBOBVoAlwcVAC8EiQCkBbEAWAVWAEoCOQCMAjX/ygRzACMIwAAaCIAAnQcAADcE4gCaBPoAAAXAAJkFxwAABcAAmwXHAJYEiQCkBbP/+gVWAJUHOwAXBQMALAXAAJkFwACZBOIAmgWdACAGqgCRBccAlgY5AFkFwACZBVYAlQXHAGEE4wAsBPoAAAbUAFkFVgAABdgAmgWfAH0ICgCaCCcAmgb1ABoH1QCdBcAAmwWxAFcIQACWBcAABARzAEkE8QBcBOsAlgNVAIgFFP/5BHMAQQWs//8D+gAYBOsAjATrAIwEAQCIBRUAGQXrAJsE1QCIBOMAUgTVAIgE4wCLBHMAVQPrABUEcwAOBwAAVARzAAwE6wCJBKUAcgarAIwGwACNBdUAKAbVAJUE6wCZBGsAOAbVAJEEq//7BHMARQTjAAADVQCIBGsAUQRzADACOQCTAkD/0AI5/6IHwAAYB0AAjATjAAAEAQCIBHMAEgTVAIgD5QCWA5MAiAgAAEEI6wCjBiAAMAAAAQEAAAAeAAAAMQAAADEAAAEBAAAAfwAAAH4AAACMAAAAjAAAAQEAAAAQAAABAQAAASEDkwB9AAAAjAJlAMgAAAMCAAD/AQKqAMkEqQBZBJsAQQOnAAoEZgAyBOoAggIvAIcDTgBaBO0AhwUDAH0CLwCHBCwAKAPtAEsD+ABBBOMAhwUKADcCLwCHAxYASwToAFAEWQAKBMAAZASyAGQD/wAKBBgACgSVAIIELAAoBbgAWgVjAC0EXgCHBF4AhwReAIcCNgBQBAkAUAaLAIcCL/+sBCwAKAQsACgD+P8WA/j/FgR5ADIFuABaBbgAWgW4AFoFuABaBKkAWQSpAFkEqQBZBJsAQQOiAAoEZgAyBOoAggKVAAADgQAABQMAfQKVAAAELAAoA+0ASwP4AEEFCgA3AxYASwToAFAEwABkBLIAZAQYAAoElQCCBCwAKAW4AFoFYwAtAi8AhwSbAEED7QBLBLIAZATbAEEAAP/cAAD/JQAA/9wAAP5RAo0AqwKNAKAC2gBDA8AAfgGW/7oAAABGAAAARgAAAEYAAABGAAAASAAAAEYAAABGAAAARgR+AYgEfgFQBH4BBAR+AJ4EfgEtBH4A6gR+ANUEfgCcBH4AvAR+AO4ENQCFAo0AwQQ1ALMGAAEABgABAAK+AFgGAAEABH4ApQR+AL0EfgDeBgABAAYAAQAGAAEABgABAAYAAQAAAABGBgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAE5v+6BgABAAYAAQAGAAEABTIAOQUyADkCLP+6Aiz/ugYAAQAGAAEABgABAAYAAQAEngA0BHgAMAQw/7oEMP+6A3YACgN2AAoGDgApBwgAKQLi/7oEVv+6Bg4AKQcIACkC4v+6BFb/ugUoAJcEbwAKA1IAAwYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAAAADAAAABGAAAARgAAAEAAAABGBgABAAYAAQAAAP/cAAD+UQAA/xYAAP8WAAD/FgAA/xYAAP8WAAD/FgAA/xYAAP8WAAD/FgAA/9wAAP8WAAD/3AAA/yAAAP/cBHMALQgAAAAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEAAo0AfwKNAGcGAAEABaAALgPAAH4B6AAAAgf/wwG8AF4B4P/6A5wABgOcAAYBvABeAeAAGgUoAJcEngARAiz/ugIs/7oBvACIAeAAGgUyADkFMgA5Aiz/ugIs/7oCvgA2A1IAAwUyADkFMgA5Aiz/ugIs/7oFMgA8BTIAPAIs/7oCLP+6BJ4ANAR4ADAEMP+6BDD/ugSeADQEeAAwBDD/ugQw/7oEngA0BHgAMAQw/7oEMP+6Ar4AaQK+AGkCvgBpAr4AaQN2AAoDdgAKA3YACgN2AAoHMgBABzIAQATe/7oE3v+6BzIAQAcyAEAE3v+6BN7/ugiAAEAIgABABiz/ugYs/7oIgABACIAAQAYs/7oGLP+6BDD/ugQw/7oEMP+6BDD/ugQw/7oEMP+6BDD/ugQw/7oEVAA0A8AARgRU/7oC4v+6BFQANAPAAEYEVP+6AuL/ugYQAC8GEAAvAnD/ugKY/7oE5gAnBOYAJwJw/7oCmP+6BFQAKQRUACkC4v+6AuL/ugOcACMDnAAjAeD/ugHg/7oC4gAhAuIAIQNS/7oDUv+6BFQAPgRUAD4CLP+6Aiz/ugK+AFgDUgADA8D/ugOc/7oDnAAGA5wABgUoAJcEbwAKBSgAlwSeABECLP+6Aiz/ugRUAAAExAAAA+QAIgRUABoD5AAiBFQAGgPkACIEVAAaBgABAAYAAQAAAABGAAAARgYAAQAGAAEABgABAAAAAEYAAABGBgABAAYAAQAAAABIAAAARgYAAQAGAAEABgABAAAAAEYAAABGAAAARgAAAEYAAABAAAAAMAYAAQAAAABGAAAARgYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAKNAMoCjQDHAo0AxgYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEAAr4AaQEA/7oIAP+6EAD/uwbTAFkFsABSBqMAkwXLAI0AAP2IAAD7wQAA/F8AAP4xAAD8rQAA/VUAAP4mAAD98QAA/RgAAPxpAAD9lQAA++AAAPxwAAD+1AAA/s0AAP6gBBsAeAasAFwGrAAZAAD+RQAA/VUAAP2mAAD8XwAA/iUAAP0YAAD74AAA+voAAPs2AAD8cAAA+4cAAPubAAD8zgAA/FQAAPvDAAD8lAAA+/UAAP2wAAD+WQAA/X4AAPyCAAD9NAAA/lAAAP5GAAD80QAA/T4AAP0CAAD8OgAA/OkAAPwmAAD8BwAA/C8AAPueAAD7dgI5AJMFxwAABHMASQXHAAAEcwBJBccAAARzAEkFxwAABHMASQXHAAAEcwBJBccAAARzAEkFxwAABHMASQXHAAAEcwBJBccAAARzAEkFxwAABHMASQXHAAAEcwBJBccAAARzAEkFVgCVBHMAQQVWAJUEcwBBBVYAlQRzAEEFVgCVBHMAQQVWAJUEcwBBBVYAlQRzAEEFVgCVBHMAQQVWAJUEcwBBAjkAagI5AF0COQCMAjkAkwY5AFkE4wBSBjkAWQTjAFIGOQBZBOMAUgY5AFkE4wBSBjkAWQTjAFIGOQBZBOMAUgY5AFkE4wBSBtMAWQWwAFIG0wBZBbAAUgbTAFkFsABSBtMAWQWwAFIG0wBZBbAAUgXHAJME4wCNBccAkwTjAI0GowCTBcsAjQajAJMFywCNBqMAkwXLAI0GowCTBcsAjQajAJMFywCNBVb//QRzAA4FVv/9BHMADgVW//0EcwAOBccAAARzAEkCOf/KAjn/ygY5AFkE4wBSBccAkwTjAI0FxwCTBOMAjQXHAJME4wCNBccAkwTjAI0FxwCTBOMAjQAA/vkAAP75AAD+9AAA/u8Eif/9A1UABwc7ABcFrP//BOIAmgQBAIgE4gCaBAEAiAXHAJYE1QCIBHMAAQRzABIEcwABBHMAEgVWAAAEcwAMBZ8AfQSlAHIFnwCcBOMAkgXPAFkEcwBMBjkAVgTjAFIFMgA5Aiz/ugJw/7oCmP+6BOYAJwIsAGUCLAAWAiwAFgIsABECLABDAiz/0gAA/vAAAAAPAAD/9QKqAJACqgCQAAAAAAAAAF4AAABeAAD/ywG8AA8B4P+/Abz/9QHg/80BvAAdAeAACQG8AIgB4AAaA5wABgOcAAYDnAAGA5wABgUoAJcEbwAKBTIAOQUyADkCLP+6Aiz/ugUyADkFMgA5Aiz/ugIs/7oFMgA5BTIAOQIs/7oCLP+6BTIAOQUyADkCLP+6Aiz/ugUyADkFMgA5Aiz/ugIs/7oFMgA5BTIAOQIs/7oCLP+6BTIAOQUyADkCLP+6Aiz/ugSeADQEeAAwBDD/ugQw/7oEngA0BHgAMAQw/7oEMP+6BJ4ANAR4ADAEMP+6BDD/ugSeADQEeAAwBDD/ugQw/7oEngA0BHgAMAQw/7oEMP+6BJ4ANAR4ADAEMP+6BDD/ugK+AE8CvgBPAr4AaQK+AGkCvgBpAr4AaQK+AE8CvgBPAr4AZgK+AGYCvgBpAr4AaQK+AGkCvgBpAr4ALwK+AC8CvgAiAr4AIgN2AAoDdgAKA3YACgN2AAoDdgAKA3YACgN2AAoDdgAKA3YACgN2AAoDdgAKA3YACgN2AAoDdgAKA3YACgN2AAoHMgBABzIAQATe/7oE3v+6BzIAQAcyAEAE3v+6BN7/ugcyAEAHMgBABN7/ugTe/7oIgABACIAAQAYs/7oGLP+6CIAAQAiAAEAGLP+6Biz/ugQw/7oEMP+6BFQANAPAAEYEVP+6AuL/ugYQAC8GEAAvBhAALwJw/7oCmP+6BhAALwYQAC8CcP+6Apj/ugYQAC8GEAAvAnD/ugKY/7oGEAAvBhAALwJw/7oCmP+6BhAALwYQAC8CcP+6Apj/ugTmACcE5gAnBOYAJwTmACcJPgAyCT4AMgdA/7oHQP+6Bg4AKQcIACkC4v+6BFb/ugRUACkEVAApAuL/ugLi/7oEVAApBFQAKQLi/7oC4v+6BFQAKQRUACkC4v+6AuL/ugYOACkHCAApAuL/ugRW/7oGDgApBwgAKQLi/7oEVv+6Bg4AKQcIACkC4v+6BFb/ugYOACkHCAApAuL/ugRW/7oGDgApBwgAKQLi/7oEVv+6A5wAIwOcACMB4P+6AeD/ugOcACMDnAAjAeD/sQHg/7EDnAAjA5wAIwHg/7oB4P+6A5wAIwOcACMB4P+6AeD/ugRUAD4EVAA+Aiz/ugIs/7oEVAA+BFQAPgRUAD4EVAA+BFQAPgRUAD4CLP+6Aiz/ugRUAD4EVAA+BJ4ANAR4ADAEMP+6BDD/ugK+AFgDUgADAxoAGgMaABoDGgAaA5wABgOcAAYDnAAGA5wABgOcAAYDnAAGA5wABgOcAAYDnAAGA5wABgOcAAYDnAAGA5wABgOcAAYDnAAGA5wABgUoAEIEb//ZBSgAlwRvAAoCLP+6Aiz/ugOcAAYDnAAGBSgAlwRvAAoCLP+6Aiz/ugUoAJcEbwAKBn8ARAZ/AEUGfwBEBn8ARQGoACgAAP4pAAD+jAAA/yUAAP8jAAD++gAA/3oAAP5ZCPwAMgitADIAAP+1AAD/tgAA/vAAAP9ZAAD+WQAA/4wBtAAAAvcAAAAA/oUAAP8HBM0AMgAA/1gAAP9YAAD/WQcyAEAHMgBABN7/ugTe/7oIgABACIAAQAYs/7oGLP+6BFQANAPAAEYEVP+6AuL/ugPAAH4C4gAhAr4AWAIs/7oCkP+6AfQALwH0ADsB9AASAfQAsQH0AG0GDgApBwgAKQIvAIcAAP7IA1AAAAReAIcD5P/1BFT/9QPkACIEVAAaA+QAIgRUABoD5AAiBFQAGgPkACIEVAAaA+QAIgRUABoD5AAiBFQAGgR+AHIEfgC9A+QADwRUAA8E4wAbBrEAHgXAAJsE4wCHBcAACgTjAAoFxwBpBccAYQRzAFUFx//9BrMAHgXAAFwE4wBUBNoATgVWAGYFAwBvBOP/rAY5AGIFGAACB3IAkgI5AJMCOQAHBccAmQRzAIkCOQAbBHMADwfvAJYFx/+tBOMAjgY5AFYHGABZBfMAVQZBAB4E4wCLBVYAlQVWAGQEcwBjBM0AWgLhAB4CqgAfBOMAGAKqAB8E4wAtBmoAYgXHAJMGKQAABHMADgTjABYEAAAiBOMAOgTjAFkENgAqBDYAOQRzADMEcwBbA/oAHgSiAB8E4wCLAj0AsAP7ALAErQBWAqoAuAqqAJQJxwCUCOMAVAlWAJ0HHACdBHIAkwo6AJgIAACYBxwAkQRzAEwFxwAABHMASQAA/v4FxwAABHMASQgA/6oHHQBYBjkAYgTjACQGOQBiBOMAVAXHAJkEcwCJBjkAWQTjAFIGOQBZBOMAUgTjADoENgAiAjn/ogqqAJQJxwCUCOMAVAY5AGIE4wBUCEMAlgVSAJUFxwCYBOMAkQXHAAAEcwBJBccAAARzAEkFVgCVBHMAQQVWAJUEcwBBAjn/NwI5/y0COf/0Ajn/5gY5AFkE4wBSBjkAWQTjAFIFxwCWAx3/zQXHAJYDHQCABccAkwTjAGcFxwCTBOMAjQVWAEoEcwAwBOMALAKqAB8EngAuBCkASQXHAJYE4wCSBZ8AnAUMAFIFDABSBOMAFgQAACIFxwAABHMASQVWAJUEcwBBBjkAWQTjAFIAAP79BjkAWQTjAFIGOQBZBOMAUgY5AFkE4wBSBVb//QRzAA4EcwBFBOMAVATjAIIE4wCHBHMANARzABQE4wBUBOMAVARzAEwGQQBMA/oATwP6ABgFhwAYBIoAUgKq/8QE4wBUBOMAVASwAFIEcwAPBM4ADwTjAIoE4wCSBOMAkgI5ABsCOQBrAz4ARAKoAAAC2QAUAjkAkwTUAJMHHQCFBx0AhQcdAH4E4/+mBOMAkQTrAIwE4wBSBqsAUgbCAE4F/wBSAx3/5gMd/+YDHf/mAx0AhwMdAIcDHQCHAx3/5gSrAIoEqwCKBHMAMAKq/8QCqv/EAqr/mwRRAB4CqgAZAqoAHwTjABsE+ABLBKgAkQRzABIGOQAJBHMADwSRAA8EAAAiBXAAIgQ2ACIENgAiBHMAQgRzAFUEcwBCBHMAVQY5AFkE6wCWBIoATwSwAFIE1QCIA6sAHgRzABQDngCIBOMAWwRzAEIEcwBVCD8AVAeJAFQJrwBUBoIAHwRGAB8GmAAfBvQAGAY1AJMFigCTBEUAHgSCAIgC8QAyAvEAMgGO/+ICBAAyAgQAAAIEAAADAAAyBC8AAALiAAAB5wBcA8sAcAI5AJgCOQB1AjkAlAKqAPMCqgDzAwAAMgMAADIErABfBKwAXwSsACoErAAqAqoBIQKqALsCqgAqAqoBIQKqABMCqgAqAqoAuwKqAMoCqgDKAqoA8wKqAPMCqgCmAqoApgKqAKYCqgATAqr/4QKq//sC7QAAASEAMgMCADIC7gAAAwAAMgMQAJYDEACWAxAAlgMQAJYDEACWAqoAYgKqAGICqgADAqoAHQQAAGkEVwCWBFcAlgRXAJYEVwCWBFcAQwRXAEMEVwBDBFcAQwRXAEMDEABDBFcALwRXAC8EVwAvBFcALwRXAC8DEAAvBFcAJQRXACUEVwAlBFcAJQRXACUDEAAvBFcAGgRXABoEVwAaBFcAGgRXABoDEAAaBFcAQgRXAEIEVwBCBFcAQgRXAEIDEABCBFcAlgRXAJYEVwCWBFcAlgRXAEIEVwBCBFcAQgRXAEIEVwBCAxAAQgRXAC8EVwAvBFcALwRXAC8EVwAvAxAALwRXAC8EVwAvBFcALwRXAC8EVwAvAxAALwRXACYEVwAmBFcAJgRXACYEVwAmAxAAJgRXAEIEVwBCBFcAQgRXAEIEVwBCAxAAQgRXAJYEVwCWBFcAlgRXAJYEVwBCBFcAQgRXAEIEVwBCBFcAQgMQAEIEVwAmBFcAJgRXACYEVwAmBFcAJgMQACYEVwAjBFcAIwRXACMEVwAjBFcAIwMQACMEVwAvBFcALwRXAC8EVwAvBFcALwMQAC8EVwBLBFcASwRXAEsEVwBLBFcASwMQAEsEVwCWBFcAlgRXAJYEVwCWBFcAQgRXAEIEVwBCBFcAQgRXAEIDEABCBFcAGgRXABoEVwAaBFcAGgRXABoDEAAaBFcAJARXACQEVwAkBFcAJARXACQDEAAkBFcALwRXAC8EVwAvBFcALwRXAC8DEAAvBFcATgRXAE4EVwBOBFcATgRXAE4DEABOBFcAlgRXAJYEVwCWBFcAlgAA/q8AAP6/AAD9tQAA/sgAAP94AAD+sQAA/z0AAP5vAAD+rgAA/84AAP9mAAD+bwAA/sgAAP7IAAD/aAAA/2gAAP9oAAAAAAAA/x8AAP8fAAD/RAAA/18AAP6HAAD/7AAA/5wAAP9RAAD/UQAA/1EAAP6/AAD/FQAAAAAAAP6xAAD/PQAA/2sAAP7yAAD/RwAA/84AAP6HAAD+uwAA/q4AAP6uAAD+yAAA/sgAAP6mAAD+vwAA/bcAAP6+AAD+pgAA/r8AAP21AAD+HwAA/uIAAP+cAAD+hwAA/0QAAP66AAD/IwAA/5oAAP25AAD+OwAAAAAAAP6nAAD/aAAA/hcAAP90AAD+hwAA/gAAAP9mAAD/RAAA/qcAAP6nAAD+pwAA/wMAAP9SAAD9HwAA/1MAAP9TAAD/UwAA/rEAAP6wAAD/oQAA/owAAP64AAD+rwAA/qIAAP66AAD99AAA/xkAAP8tAAD+jAAA/ogCqgC7AqoAKgKqAMgE4gBnBKgACgYpAAAIAgAABikAAAX/AFIGwgBOBWkAFAY5AFkE4wBSBccAdwRzAFUE4wCXA54AiAYDAAAEPAAdBm8ACgTiAAoH7wCWBx0AhQWfAH0E4wCKBZ8AnATXAAoFVgBkBVYAZAUkABQE1AAKBeEAVQSgAEsEDgAUA4QAKAVpABQE8QBcBHMAVQI5/6IGOQBWA9QAUQPUAFEFVgCVBcAAmQRzAEEE6wCMCj0AWQY6ABQG9AAaBZ8AGwfOAIwGXgCTBVYAAARzAAsHaACMBmcAkwZ5AFYGBwB2CJ4AjAfYAJMFAwBGA/oAQwZ5AFYGBwB2BjkAVgTjAFIGhf//BSwACwaF//8FLAALCPYAWQfLAFIGhAAjBRoAIwo9AFkHNQBVAAD+Nwo9AFkGOgAUBccAYQRzAFUErAAPAAD+pgAA/rEAAP+NAAD/jQAA/CsAAPxMBcAAmQTrAIwFwAARBOsAGwVWAJUE4wCLBZ8AnATJAIgFAwAsA/oAGATiABEEAQANBhcAGgT8ACgHCQCWBbYAiAkCAJkHXwCIBccAOwSfADQFxwBhBHMAVQTjAC0D6wAVBtIALAWDABUFnwB9BKUAcgbaAAoFbQAKBtoACgVtAAoCOQCMBzsAFwWs//8FnQCaBMgAiAWdACAFFQAZBccAlgTVAIgFxwCWBNUAiAWfAH0EpQByBqoAkQXrAJsCqgAaBccAAARzAEkFxwAABHMASQgA/6oHHQBYBVYAlQRzAEEFzwBZBHMATAc7ABcFrP//BQMALAP6ABgFAwAsBDYAIgXAAJkE6wCMBcAAmQTrAIwGOQBZBOMAUgY5AFYE4wBSBbEAVwRrADgE+gAABHMADgT6AAAEcwAOBPoAAARzAA4FnwB9BKUAcgfVAJ0G1QCVBcAAXgTjAFQIPgBeB3oAVAetAEYGxABDBUMARgRKAEMIGgAgB6UAGQhDAJYHZgCIBjkAYgSwAFIGIAAtBZsAFQAA/0MAAP7JAAD/dwAA/7AAAP9HAAD/VgAA/3QAAP7XAAD+rAAAAAAAAP9SAAD/VgAAAAAAAP6sAAD9mgAAAAAAAP9qAAD/fAAA/2kAAP9WAAD+rAAA/38AAP9WAAD97wAA/0MAAP9pAAD/fAAAAAAAAP2uAAD/jAAAAQIAAP7vAAD+7wAA/v0AAP75AAD/UwAA/vgAAP75BccAAARzAEkFxwCWBOMAhwXHAJYE4wCHBccAlgTjAIcFxwBhBHMAVQXHAJQE4wBUBccAlATjAFQFxwCUBOMAVAXHAJQE4wBUBccAlATjAFQFVgCVBHMAQQVWAJUEcwBBBVYAlQRzAEEFVgCVBHMAQQVWAJUEcwBBBOMAlwKqABgGOQBiBOMAVAXHAJYE4wCSBccAlgTjAJIFxwCWBOMAkgXHAE4E4wA7BccAlgTjAJICOf/SAjn/0gI5ABsCOf/OBccAmQRzAIkFxwCZBHMAiQXHAJkEcwCJBOMAnQI5AJME4wCdAjn/6wTjAJ0COf/dBOMAnQI5/8sGqgCRBx0AfgaqAJEHHQB+BqoAkQcdAH4FxwCYBOMAkQXHAJgE4wCRBccAmATjAJEFxwCYBOMAkQY5AFkE4wBSBjkAWQTjAFIGOQBZBOMAUgY5AFkE4wBSBVYAlQTjAIsFVgCVBOMAiwXHAJYDHQCHBccAlgMdAIcFxwCWAx0AhwXHAJYDHQBZBVYASgRzADAFVgBKBHMAMAVWAEoEcwAwBVYASgRzADAFVgBKBHMAMATjACwCqgAfBOMALAKqAB8E4wAsAqoAHwTjACwCqgAfBccAkwTjAI0FxwCTBOMAjQXHAJME4wCNBccAkwTjAI0FxwCTBOMAjQVW//8EcwALBVb//wRzAAsHjQAHBjkACQeNAAcGOQAJBVYAAARzAAwFVgAABHMADAVW//0EcwAOBOMAFgQAACIE4wAWBAAAIgTjABYEAAAiBOMAkgKq/94GOQAJBHMADgRzAEkCOQCNBOsATgTrAE4E6wBOBOsATgTrAE4E6wBOBOsATgTrAE4FxwAABccAAAbz//IG8wAABvP/8gbzAAAG8wBDBvMAQwPMAE4DzABOA8wATgPMAE4DzABOA8wATgYe//IGHgAAB67/8geuAAAHrv/yB64AAATjAI4E4wCOBOMAjgTjAI4E4wCOBOMAjgTjAI4E4wCOBo//8gaPAAAIH//yCB8AAAgf//IIHwAACB8AFAgfABQCOQCQAjkAkAI5/7YCOf/EAjn/3gI5/+wCOf+zAjn/wAMB//IDAQAABJH/8gSRAAAEkf/yBJEAAASRABQEkQAUBOMAUgTjAFIE4wBSBOMAUgTjAFIE4wBSBp3/8gadAAAIVf/yCFUAAAfJ//IHyQAABKgAdgSoAHYEqAB2BKgAdgSoAHYEqAB2BKgAdgSoAHYGggAAB/4AAAhiAAAHrv/zBsIATgbCAE4GwgBOBsIATgbCAE4GwgBOBsIATgbCAE4Gzv/yBs4AAAiG//IIhgAAB/r/8gf6AAAH+v/zB/r/8wTrAE4E6wBOA8wATgPMAE4E4wCOBOMAjgI5/+cCOQCNBOMAUgTjAFIEqAB2BKgAdgbCAE4GwgBOBOsATgTrAE4E6wBOBOsATgTrAE4E6wBOBOsATgTrAE4FxwAABccAAAbz//IG8wAABvP/8gbzAAAG8wBDBvMAQwTjAIwE4wCMBOMAjATjAIwE4wCMBOMAjATjAIwE4wCMBo//8gaPAAAIH//yCB8AAAgf//IIHwAACB//8wgf//MGwgBOBsIATgbCAE4GwgBOBsIATgbCAE4GwgBOBsIATgbO//IGzgAACIb/8giGAAAH+v/yB/oAAAf6//MH+v/zBOsATgTrAE4E6wBOBOsATgTrAE4E6wBOBOsATgXHAAAFxwAABcf/0QXH/90FxwAAAqoA3AKqAMoCqgDcAqr/8wKq//ME4wCMBOMAjATjAIwE4wCOBOMAjAbmAAAG5gAAB1cAAAdXAAAFxwCWAqr/8gKq//ICqv/zAjn/5QI5/9sCOf/OAjn/zgI5/8ICOf+7Ajn/6AI5/94DyQAAA8kAAAKqAAACqgAAAqr/8wSoAHYEqAB2BKgAdgSoAHYE8wB2BPMAdgSoAHYEqAB2BVb//QVW//0G5v/YB0r/3QYeAAADuP/0A7j/9AKqACoGwgBOBsIATgbCAE4GwgBOBsIATgdl/9EGnf/dB5b/0QbO/90GagBiAqoAuwKqANwEcwAKBccAYQXHAGEHHQB+BccAIQnNAJYHjQAHBccAIATjAC0IsAAUBAAAMATBAGYAAP9TAAD/UwAA/1MAAP9TAjkAGwI5/6IEcwAABVYAEgazAFQD/gBXBqsAkQQMAB8F1v/mBdb/5gKqAIQCqgCEAqoAyQKqAMkCqgCRAqoAKgKq/8UCqv/DAqr/8wKqAMkCqgCpAqoAqQKqAKkCqgCpAy4AHgMuAB4CqgA6AAD/cwAA/50AAP7IAAD/IwAA/3IAAP9yAAD+5wAA/50AAP9TAAD/UwAA/1MFVgCVBOMAiwS1AAAGNQAABx0AYQTrAA8EcwBVBJkAkQSZABsEAQCMA/oAGAI5AJMEDwBJBHYAjgOeAA4F6wCbBOsAjATjAFIEcwA0BPEAUgTxAFIE8QAhB40AVASSAEsE4wBTBOMAUwTpAIwEq//7BKv/+wPrABUEqAB2BOMAUQYkAFEE4ABRBHMACwY5AAkEAAAiA98AIgPyAEsE7AAUA1UAiARzABIE1QCIBOkAjAYHAHYFFQAZA+MAAAWRAAADogAyA6IAAAOjADIDVQAyA1UAMgQDADIDfAAyAXIAVQLeADIDsAAyAx4AMgQiADIDdwAyA3gAMgQmADIDegAyA1sAMgOsADIDdwAyA3sAMgUUAAADBQAyAwUAMgMhADIEtgAyAyEAMgMhADIDAgAyAwIAMgLPADICzwAyAyAAMgEhADICygAyBIQANALyADIDSAAyAwoAMgNJADIDSQAyAyAAMgG8AAoC8gAyA0IAMgSEADIC6QAAA0wACgMbADIC6QAAA0MAMgPaADIDCAAAASEAMgIEADIC8gAyAukAAAMbADIC6QAAA0IAMgPaADIDCAAABe0ARgqYAEYGEwBGBon/ugVB/7oB6QAeBFQAEAAA/w0AAP81AAD+zgAA/rcAAP7JAAD/xwAA/08AAP+eAAD+8AK+AGkCvgBpA3YACgN2AAoDwP+6A5z/ugPA/7oDnP+6BcgAOQWSADIGFgCCBRkASwUkAEEGDwCHBVgAKAaPAC0ErABVAAD+OwAA/mYAAP5oBHP//AQAAIQD1f+6AeD/ugHg/7EB4P+6AeD/ugbQAC4JhAAjBAAAAAgAAAAEAAAACAAAAAKrAAACAAAAAVUAAARzAAACOQAAAZoAAACrAAAAAAAABeX/9wXHAGEGqgCRBesAmwdgAI0HoQBUB6EAWwXHAAAFxwBhBHMAFATjABEE4wAsBHMAOQQAACIFKQBCAAABAQAA/0IAAP6tAAD/OgAA/1ME8wAKBccAaQXHAGEFxwBpBIkApANVAIgAAP9DAAD/AQAA/6wDFgB9AAD/NwKY/7oDPQAeAAD/OgAA/0gAAP9JAAD/fgAA/08AAP9KAAD+ngUyADkFMgA5Aiz/tgIs/7YFMgA8BTIAPAIs/7oCLP+6BTIAOQUyADkCLP+6Aiz/ugUyADkFMgA5Aiz/ugIs/7oFMgA5BTIAOQIs/7oCLP+6BTIAOQUyADkCLP+6Aiz/ugUyADkFMgA5Aiz/ugIs/7oEngA0BHgAMAQw/7oEMP+6BJ4ANAR4ADAEMP+6BDD/ugK+AE8CvgBPAr4AaQK+AGkDdgAKA3YACgcyAEAHMgBABN7/ugTe/7oEVAA0A8AARgRU/7oC4v+6BFQANAPAAEYEVP+6AuL/ugRUADQDwABGBFT/ugLi/7oGEAAvBhAALwJw/7oCmP+6BhAALwYQAC8CcP+6Apj/ugYOACkHCAApAuL/ugRW/7oGDgApBwgAKQLi/7oEVv+6Bg4AKQcIACkC4v+6BFb/ugLiACEC4gAhA1L/ugNS/7oC4gAhAuIAIQNS/7oDUv+6BFQAPgRUAD4CLP+6Aiz/ugRUAD4EVAA+Aiz/ugIs/7oEVAA+BFQAPgIs/7oCLP+6A5wAIwOcACMB4P+6AeD/ugN2AAoDdgAKA3YACgN2AAoHMgBABzIAQATe/7oE3v+6BOP/wQTjAFQCqv/zBx3/wQTj/9UE4//FAx3/wQMd/8EEc///Aqr/2gQAACEE4wCDAvAAMgTcAE4G+wAfAjkAGwI5ABsE4wAUBKgAFAT4ABQE4wCHBOMAVAKqABgGJQBUBHMAiQI5AHAHHQB+BOMAkQTjAIsDHQBmBHMAMAO6/8QEcwALBHMADAQAACIEcwBJBOMAVATjAFQEcwBBA/oATwP6ABgFPgBRAjkAkwRzADQCqv/EBOMAjQQ2ACIDIQAyAwoAMgMKAAYDSAAyAs8AMgHwAAoB8AAAAyAAMgLxADIBdAAKASEAMgEhADIBdAAKAnYAAAGOADIBUAAyAkkAMgSEADQEhAAyA18AAANfADIC+gAyA0gAMgQDADIDAgAyAjkAAAG8AAoDQAAKA14AMgLqADIC6gAyAukAAALkADIC5AAyA74AMgMKADIC6AAyAAD+kgAA/pIAAP9zAAD+nwKqAMkDBQAyAwIAMgNIADIC7gAAAwIAMgY5AGIFxwAABVYAHgXHAGECqgBBBOsATgTrAE4E6wBOBOsATgTrAE4E6wBOBOsATgTrAE4COf+2Ajn/tgI5/8QCOf/EAjn/tgI5/7YCOf/EAjn/xASoAHYEqAB2BKgAdgSoAHYEqAB2BKgAdgSoAHYEqAB2Ajn/yQI5/8kCOf/JAjn/yQSoAHYEqAB2BKgAdgSoAHYD5AAiBFQAGgPfADAFx//9BccAFgVWAAAFVgCVBHMAQQRzACMCOf+iBjMAWQTjAFsFxwAAAx0AGwVW//0EcwAOBHMANARzAFUEcwA0AjkAkwSJABEDVQAbBVYAAARzAAwFVgAABHMADAUDAG8D+gBPBZ0AIAUVABkAAP7GAAD+1AAA/sYAAP7UAAD+XwAA/l8AAP9yAAD/cwAA/ucIAAAABAEAXQRzADQE4wARAjkAGwTjAAYFVv/9BccAlgRzAEkCqv/NBccAlgTjAJIFxwCZBHMAiQTjABYEAAAiBHMAKARUAJYDfACIBbkATgAA/1MAAP+8AAD+/gAA/v4AAP6kAAD+pAI5AJMFyQCcBccAmAXJAJwAAP7gAAD/MAAA/tQAAP7VAAD+wAAA/tAAAP7YAAD+2AAA/tgAAP7YAAD9xgY5AFkE4wBbB40ABwY5AAkFuQCRAAD+mwYbAFkE2QAGCFsABwbeAAYCqgDJAxwAVQHnAFwB5wBcBAAAmQQAAJkCqgC4AqoAuAKqALgCqgADBOMALARzACsEwwAKBHMAFAaXAIcHOABQAAAAAAAAAGwAAABsAAAAbAAAAGwAAABsAAAAbAAAAGwAAABsAAAAbAAAAGwAAABsAAAA9gAAAYAAAAGAAAABgAAAAYAAAAGAAAABvgAAAhQAAAMYAAADmgAABUAAAAaYAAAHsgAACSQAAApYAAALFAAADLIAAA34AAAN+AAADfgAAA34AAAN+AAADfgAAA34AAAN+AAAD3IAABDaAAASFAAAEv4AABO8AAAUWAAAFZ4AABZyAAAW+gAAFvoAABjEAAAZIAAAG3QAAB1yAAAeegAAH0oAAB9KAAAgrgAAIw4AACOkAAAkhAAAJIQAACSEAAAkhAAAJXoAACV6AAAl7gAAJe4AACXuAAAl7gAAJe4AACXuAAAn/AAAKPgAACo0AAArJAAALTAAAC4wAAAwDAAAMQwAADGuAAAxrgAAMa4AADIaAAAzzgAANLgAADWoAAA2pAAANqQAADeIAAA6zgAAO+4AADzWAAA+KgAAQEYAAEIcAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAEOaAABDmgAAQ5oAAQAADV0A8gA8AI8ABgACABAALwBVAAAHPP//AAUAAgAAABQA9gABAAAAAAAAABAAAAABAAAAAAABABEAEAABAAAAAAACAAcAIQABAAAAAAADABEAKAABAAAAAAAEABEAOQABAAAAAAAFAAwASgABAAAAAAAGABEAVgABAAAAAAAHAAcAZwABAAAAAAAIAAcAbgABAAAAAAAJAAcAdQADAAEECQAAACAAfAADAAEECQABACIAnAADAAEECQACAA4AvgADAAEECQADACIAzAADAAEECQAEACIA7gADAAEECQAFABgBEAADAAEECQAGACIBKAADAAEECQAHAA4BSgADAAEECQAIAA4BWAADAAEECQAJAA4BZk9yaWdpbmFsIGxpY2VuY2VCT0dBSkMrQXJpYWwsQm9sZFVua25vd25CT0dBSkMrQXJpYWwsQm9sZEJPR0FKQytBcmlhbCxCb2xkVmVyc2lvbiAwLjExQk9HQUpDK0FyaWFsLEJvbGRVbmtub3duVW5rbm93blVua25vd24ATwByAGkAZwBpAG4AYQBsACAAbABpAGMAZQBuAGMAZQBCAE8ARwBBAEoAQwArAEEAcgBpAGEAbAAsAEIAbwBsAGQAUgBlAGcAdQBsAGEAcgBCAE8ARwBBAEoAQwArAEEAcgBpAGEAbAAsAEIAbwBsAGQAQgBPAEcAQQBKAEMAKwBBAHIAaQBhAGwALABCAG8AbABkAFYAZQByAHMAaQBvAG4AIAAwAC4AMQAxAEIATwBHAEEASgBDACsAQQByAGkAYQBsACwAQgBvAGwAZABVAG4AawBuAG8AdwBuAFUAbgBrAG4AbwB3AG4AVQBuAGsAbgBvAHcAbgAAAAMAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAACxVIBBDQOsAK8DrAACABADrAAgA6wAoAOsAAMAQAOsswcNMkC4A6yzEhQyQLgDrLIWKzK5/8ADrLI6M0C4A6yzLZQygLwDqwBfADP/wAOrslUzQLgDq7NARDJAuAOrszM7MkC4A6uzLzEyQLgDq7IIM0C4A6uzBxQyH0EaA6sALwOrAAIADwOrAC8DqwBPA6sAjwOrAJ8DqwC/A6sABgAQA6sA3wOrAP8DqwADA6gDorJGH0C4A6WyCDMPQRQDpQABAEADpQDPA6UA/wOlAAMAIAOlAK8DpQDvA6UA/wOlAAT/wAOjswkMMkC4A6OyCDMPQRsDowABAA8DowAQA6MAgAOjAK8DowDPA6MABQBvA6MAnwOjAP8DowADAJ8DogCvA6IAAgOiA6GyEB8QQQoDngB/A54AAgOaAA8BAQAf/8ADmLMQFDJAuAOZsw8TMkBBEAOVAFADlQACALADTQDAA00AAgBvA5EAfwORAAL/wANLsi0xMrn/wANLswoOMhBBEAOLACADiwCAA4sAAwCgA4sAAQAgA4sAQAOLAAL/wAOLsxMWMkC4A4OyDxEyuf/AA3uyMDQyuf/AA3uzEBgyUEEUA3gAAQNlA24AIwAfA34DbgAeAB8DYwNuAB0AHwNiA2QADQAf/8ADQLMPEDKAQRADPwABAz8DFQApAB8DQQMWADIAHwNEAxoAGwAf/8ADdbIOETK5/8ADdbIoKjJBCgNDAxgAMgAfAw8DDQA0AB8DCAMHsjIfILsDQAABAEADiLMJCzJAuAOIshAVMr0DhQMHABQAHwOAAweyFx8PvQMKAC8DCgAC/8ADVLMJDTKQQQwDVACgA1QAAgAfA24AAQCfA24AAQBAA26yCQsyQREDRQMcABYAHwNrAx0AFQAfA0YDHgAVAB8DpwOhAEYAHwOdsyYcH8C7A5MAAQBAA5KzCQ0yQLgDPrIIM0C4Az6zDQ4ywEEJAz4AAQCwA44AwAOOAAL/wAOQsyY4MgBBJgMoADADKAACACADfwAwA38AAgAQA4oAMAOKAFADigBvA4oAfwOKAJ8DigAGAAADiQAwA4kAAgAvA3oAcAN3AJADdwCfA3oABP/AAxWyDxAyuf/AAxWyJCgyuQMZAxiyMh8QuwMaAAH/wAMaswkOMkC4AxiyEhMyuf/AAxizDA4yP70DcwBPA3MAAgBAA3SzFxgyb7sDKgABAEADLLMYGzJAuANwsgkMMr0DFwMWADIAH//AAxayDhEyvQMcAx4AFgAfAx0DHrIVH7BBHwMeAAEADwMfAAECygLQABUAHwLTAtUADQAfAs8C0AANAB8CywLQAA0AHwLNAtAADQAfAs4C0AANAB//wALQswkMMkC4AtKzCQwy4EEcAuUAAQBfAt0AnwLlAAICuwLDADAAHwLaArgAMgAfAtkCuQA/AB8C2AK4AGQAHwK5ArgAMwAfArqyIcgfuAK4syHIH0C4A5uyDRYyuf/AAsOyKy8yuf/AAsOyHyUyuf/AAsOyFxsyuf/AAsOyEhYyQSUCwgLBABwAHwLXAsEAJAAfAsECwAAiAB8CvwLAABgAHwLAAnQAyAAfArUCNQA7AB8CtAI1ADsAHwLEArwAHgAfArcCtgA4AB8Cs7IOyB+4ArCyB8gfuAKvsgbIH7gCrrIAyB+4Aq+yUC8fvAKuAqsAGgAfAq2yJhofuAKosyYkHw+7AjUAAQKlAnSyHR8SQQoCoQFYAfQAHwKgANgB9AAfABICorI3yB+4ApCyvCAfuQKQApBAGDdAJUAtQKYDMCUwLTCmAyAlIC0gNyCmIEEQAo4ABQCfAosAAQKLAosANwAgAokAMAKJAEACiQCQAomyBDewQf0CdADAAnQAAgCAAnQAoAJ0AAIAYAJ0AHACdAACAAACdAAQAnQAAgCAAnQA8AJ0AAIAPwKFAE8ChQACAJACfgCQAn8AkAKAAJACgQAEAJACegCQAnsAkAJ8AJACfQAEAJACdACQAnUAkAJ3AAMAcAJ+AHACfwBwAoAAcAKBAAQAcAJ6AHACewBwAnwAcAJ9AAQAcAJ0AHACdQBwAncAAwBgAn4AYAJ/AGACgABgAoEABABgAnoAYAJ7AGACfABgAn0ABABgAnQAYAJ1AGACdwADAFACfgBQAn8AUAKAAFACgQAEAFACegBQAnsAUAJ8AFACfQAEAFACdABQAnUAUAJ3AAMAQAJ+AEACfwBAAoAAQAKBAAQAQAJ6AEACewBAAnwAQAJ9AAQAQAJ0AEACdQBAAncAAwAwAn4AMAJ/ADACgAAwAoEABAAwAnoAMAJ7ADACfAAwAn0ABAAwAnQAMAJ1ADACdwADACACfgAgAn8AIAKAACACgQAEACACegAgAnsAIAJ8ACACfQAEACACdAAgAnUAIAJ3AAMAEAJ+ABACfwAQAoAAEAKBAAQAEAJ6ABACewAQAnwAEAJ9AAQAEAJ0ABACdQAQAncAAwDgAn4A4AJ/AOACgADgAoEABADgAnoA4AJ7AOACfADgAn0ABADgAnQA4AJ1AOACd7ED0EHFAn4A0AJ/ANACgADQAoEABADQAnoA0AJ7ANACfADQAn0ABADQAnQA0AJ1ANACdwADADACdABAAnQAAgDAAn4AwAJ/AMACgADAAoEABADAAnoAwAJ7AMACfADAAn0ABADAAnQAwAJ1AMACdwADALACfgCwAn8AsAKAALACgQAEALACegCwAnsAsAJ8ALACfQAEALACdACwAnUAsAJ3AAMAoAJ+AKACfwCgAoAAoAKBAAQAoAJ6AKACewCgAnwAoAJ9AAQAoAJ0AKACdQCgAncAAwCQAn4AkAJ/AJACgACQAoEABACQAnoAkAJ7AJACfACQAn0ABACQAnQAkAJ1AJACdwADACACfgAgAn8AIAKAACACgQAEACACegAgAnsAIAJ8ACACfQAEACACdAAgAnUAIAJ3AAMCgQFYCAEAHwKAASkIAQAfAn8A7AgBAB8CfgDYCAEAHwJ9ALEIAQAfAnwApggBAB8CewCCCAEAHwJ6ADcIAQAfAncAJggBAB8CdQAgCAEAHwJ0AB8IAbIfNw9BFgI1AE8CNQBfAjUAbwI1AJ8CNQCvAjUAvwI1AAcArwI1AM8CNQDfAjUA/wI1QCIEDwdPB58Hrwe/BwWvB+AHAg8GTwafBq8GvwYFrwbgBgIgQRsCDQABAF8CNQABAI8CNQABAH8CNQDvAjUAAgAvAjUAPwI1AAIAPwI0AE8CNAACAjUCNQI0AjRAEe0g7yoBzyoBvyoBryoBjyoBQQkCRwEEAB4AHwIgADcCAQAfAVhADCY+H9gmPh83Jic+H7gCjrbsFx+yJjYfuAG8siY2H7gBKUArJjYf7CY2H7EmNh+mJjYfgiY2HzcmNh8yJjYfLSY2HyUmNh8fJjYfNyYqH7gBWEAiJj4f2CY+H7wmPh8nJj4fISY+HyAmPh83ABYWAAAAEhEIQLkCDQGms8UNAAm4AbyyJygfuAG7sicwH7gBuLInTx+4AbeyJ2IfQQkBtgAnAQEAHwG1ACACqwAfAa+yH+QfuAGtsh/kH7gBrLIfux+4AaiyHzQfuAFdsicuH7gBW7InzR9BDQFVAB8EAQAfAVQAHwQBAB8BUwAfAgEAHwFSsh9WH7gBUbIfKR+4ASuyJyYfQQ0BKgAnASUAHwEpAVgA5AAfASUAHwQBAB8BJLIf5B+4ASOyHzsfuAEish85H0ENAQgAJwgBAB8BBgAtAQEAHwEFAB8BAQAfAQOzH7sf77kBWAQBQAsf7R+TH+wf5B/rH7gCAbIf2SC4BAGyH88luAFWQAofvC2eH7sfQR+yQQoBWAQBAB8AsQFYBAEAHwCwAVgEAbUfpiWJH5u5AVgBJbYfmR8uH44tuAgBtR+NHykfibkBWAQBsh+CILgCq0ATH4AfMB90LeQfcx9KH2EfUh9dJbgCq7IfXB+8CAEAHwBZAVgCq7YfUCWJH0kfuAElsh9HJbgEAUALH0YfeR9AHycfOSC8AqsAHwA4AVgEAbIfNy28ASUAHwAyAVgBJbYfLB80HyoluAgBsh9VN7gBEUAqB/AHkAdbB0IHOwcjByIHHgcdBxQIEggQCA4IDAgKCAgIBggECAIIAAgUuP/gQCsAAAEAFAYQAAABAAYEAAABAAQQAAABABACAAABAAIAAAABAAACAQgCAEoAsBMDSwJLU0IBS7DAYwBLYiCw9lMjuAEKUVqwBSNCAbASSwBLVEKwOCtLuAf/UrA3K0uwB1BbWLEBAY5ZsDgrsAKIuAEAVFi4Af+xAQGOhRuwEkNYsQEAhY0buQABARmFjVlZABgWdj8YPxI+ETlGRD4ROUZEPhE5RkQ+ETlGRD4ROUZgRD4ROUZgRCsrKysrKysrKysrGCsrKysrKysrKysYKx2wlktTWLCqHVmwMktTWLD/HVlLsIFTIFxYuQIPAg1FRLkCDgINRURZWLkEcAIPRVJYuQIPBHBEWVlLsORTIFxYuQAgAg5FRLkAJwIORURZWLkIQgAgRVJYuQAgCEJEWVlLuAElUyBcWLkAJgIPRUS5ACECD0VEWVi5Cg0AJkVSWLkAJgoNRFlZS7gEAVMgXFix2CBFRLEgIEVEWVi5JQAA2EVSWLkA2CUARFlZS7gEAVMgXFi5AVgAJkVEsSYmRURZWLkjIAFYRVJYuQFYIyBEWVlLsClTIFxYsR8fRUSxLR9FRFlYuQENAB9FUli5AB8BDURZWUuwL1MgXFixHx9FRLElH0VEWVi5ATUAH0VSWLkAHwE1RFlZS7gDAVMgXFixHx9FRLEfH0VEWVi5FCgAH0VSWLkAHxQoRFlZKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrK2VCKwGzMXV+w0VlI0VgI0VlYCNFYLCLdmgYsIBiICCxfnVFZSNFILADJmBiY2ggsAMmYWWwdSNlRLB+I0QgsTHDRWUjRSCwAyZgYmNoILADJmFlsMMjZUSwMSNEsQDDRVRYscNAZUSyMUAxRSNhRFmzPzxYQUVlI0VgI0VlYCNFYLCJdmgYsIBiICCxWDxFZSNFILADJmBiY2ggsAMmYWWwPCNlRLBYI0QgsT9BRWUjRSCwAyZgYmNoILADJmFlsEEjZUSwPyNEsQBBRVRYsUFAZUSyP0A/RSNhRFlFaVNCAUtQWLEIAEJZQ1xYsQgAQlmzAgsKEkNYYBshWUIWEHA+sBJDWLk7IRh+G7oEAAGoAAsrWbAMI0KwDSNCsBJDWLktQS1BG7oEAAQAAAsrWbAOI0KwDyNCsBJDWLkYfjshG7oBqAQAAAsrWbAQI0KwESNCACsrKysrKysrALASQ1hLsDVRS7AhU1pYsSYmRbBAYURZWSsrKysrKysrKysrKysrKysrKytzc3Nzc0WwQGFEGABFaURFaURzc3N0c3NzdHN0c3QrKysrKysrKysrKysAc3Nzc3Nzc3Nzc3Nzc3Nzc3Nzc3Nzc3R0dHR0dHR0dHR0dHR0dHR0dHR0dHV1dXN0dXV1dStzAABLsCpTS7A2UVpYsQcHRbBAYERZAEuwLlNLsDZRWlixAwNFsEBgRLEJCUW4/8BgRFkrRWlEAXQAc3NzK0VpRCsBK0NcWEAKAAYABwKgBqAHArn/wAJ0sxodMm+9AncAfwJ3AAL/wAJ3si8xMrn/wAJ3syIlMkC4AnSzLzUyQLgCdLMoKjJAuAJ0shohMrj/wLM3Gh0yuP/AsyUaHTK4/8BAES0aHTKQJZAtkDegJaAtoDcGuP/AtqYaHTIfph+4Ao6yL6YDAHQrcysrKysrKysrdCtzdFkAKytDXFi5/8ACobIcHTK5/8ACoLIcHTIrK1krcwErKysrACsrKysrKysrKysrKysrKysrKwErKysrKysrc3QrKysrKysrK3NzKysrKysrcytzKysrdCsrK3Nzc3NzK3NzKysrcysrACsrKytzdHMrcysrKyt1KysrKysrKyt1KysrKytzKysrK3N0dSsrc3NzKysrcytzc3R1KytzdHUrK3N0dSsrKysrKysrKysrK3R1KwAA); }&#xA;@font-face { font-family: &quot;g_font_2&quot;; src: url(data:font/opentype;base64,AAEAAAANAIAAAwBQT1MvMmJoWKEAAADcAAAATmNtYXCkFUN4AAABLAAAAJhjdnQgoRzX6wAAAcQAAAZUZnBnbcx5WZoAAAgYAAAGbmdseWYy9I76AAAOiAAAb2hoZWFk53kpCAAAffAAAAA2aGhlYRIzFiYAAH4oAAAAJGhtdHh0wP1UAAB+TAAANXRsb2NhBbbUQAAAs8AAADV4bWF4cBK5AcEAAOk4AAAAIG5hbWUOcFvzAADpWAAAAi5wb3N0AAMAAAAA64gAAAAgcHJlcCXWTb8AAOuoAAALvgAABAABkAAFAAAEAAQAAAAEAAQABAAAAAQAAGYCEgAAAQEBAQEBAQEBAQAAAAAAAAAAAAAAAAAAAAA/Pz8/AEAAIACpCAACAADMCAwDmAAAAAAAAQADAAEAAAAMAAQAjAAAAB4AEAADAA4AIAAlACkAOgA9AD8ASQBaAF8AaQB6AKkgE+AB//8AAAAgACUAKAArAD0APwBBAEwAXwBhAGsAqSAT4AD////j/+P/4//j/+P/4//j/+P/4//j/+P/4uCeAAAAAQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAQAAAADABAFugAZBboAGgWnABkEJgAYAAD/5wAA/+gAAP/n/mn/6AW6ABn+af/oAuoAAAC4AAAAuAAAAAAAqACtAWkArQC/AMIB8AAYAK8AuQC0AMgAFwBEAJwAfACUAIcABgBaAMgAiQBSAFIABQBEAJQBGf+0AC8AoQADAKEAzQAXAFcAfgC6ABYBGP/pAH8AhQPTAIcAhQANACIAQQBQAG8AjQFM/3UAXADfBIMANwBMAG4AcAGA/1j/jv+S/6QApQC5A8j//QALABoAYwBjAM3/7gXY/9wALQBcAJUAmQDfAZIJtQBAAFcAgAC5A50AcgCaA10EAf9n//oAAwAhAHcAzQAEAE0AzQHAAisATABlAOcBGAF8A0MF2P+j/7D/xAADABwAXQBoAJoAugE1AUcCIQVc/03/zQAWAC0AeACAAJkAsgC2ALYAuAC9ANoBDAXw/6T/8AAZACwASQB/ALQAzgHAA/79gf4/AAAABQAYACkAOQBJAG8AvgDHANABIwHBAm8FDAUyBUAFev/UABQAMQBVAFcApwC0AOYB9wJ+An4CfwPGBEb/QgAOAIUAkQC/AMIAxQDhARoBLwFPAVYCKQJvAp4DcgAIACwAMQAxAGQAaQCJAJgAxwDeASsBtgIMAs8DowSrBPsGHf7g/w4ABgAmAJsAnQDBAQ0BGAEgAXMBggHWAeMCQwJfApsC4gOUBKkE0gdhABwAXgBtAI0AqwD3ARIBOAFRAVsBaAF8AYcBkQGZAc0B0AHoAkECVAJrAu8DaANxA70EQgRCBFMEcwSDBYYFiwbo/lj+xP7R/vf/Mv+GAFEAfACBAJEAlQCeALQAuQDPANkA2QDfAOIBBQELAQ4BDgEgASEBVQF7AXsBfgGNAaIBqAGpAbQB0AHQAeIB6QHyAfUB+wIAAgACBgIbAiECIgIiAiMCcgJ3ApQCnALPAs8C0ALsAvkDFwMiAysDNQM8A1kDbwNxA4cDkAOQA7UD4QQaBM8E/wUyBTIFlgWfBagFqwXCBfAGDAeCCAAIzPyj/Sr93v4A/oj+lv6y/rT/4QAVABkAGgAcAB8APABRAGEAYQBqAHgAlgClAK8A0wEMARgBGgEqAT4BTAFRAV8BagFxAXgBggGEAZoBpQGoAakBrgG8Ac0B1wHvAgACDQIcAiECIgIuAjUCQgJPAk8CXgJlAnECkAKSArQC1gL6AwcDCwMPAxUDKgNHA10DZQN0A3kDlgOwA8wD3QPiA/YD/AP8A/8ECgQfBCIEJgQrBEcEXwR1BJ4E5wTnBVwFywXlBgoGbQaGBrgG8Qc2Bz4HUAdRB10Hjwe2B9QIYAC2AMMAtQC3AAAAAAAAAAAAAAAAAeADgQNFA7UAjgIzBBkCzgLOAC0AXwBkA00CPwAAAqgBiAJ9AbQCJAV4BjsCOwFOAPAEJgKUAsYCnwL2AjsDTQFLAVMAagIxAAAAAAAABhQEqgAAADwEwwDtBLwCZQLOA7UAeAYMAX4C7wYMALIBAAI5AAABxQMwBCsDywDaA98BBwShANsECgEXAe0CpwNQAQsBvQQ+BVgAIQOcAK4DcQF9ALUCRQAACvsIjAErAU4BqgCHAFQBMgH4A/8AAwJOALQANwPjAIMAawLYAO0AdwCIAJcBZARnAI4AMwF8AOcApgKeAykFbgYqBhUByQJpBIoCEwG0AAIEqQAAAjkBJAEDBRQAhAFdA5oG7wLZAHUAzwQKAN4DrAS8As8CrgNNBPAFUgFoAG0AfQCGAHH/gQB5BVgE0gFnAAMBVgAlBOAAlAB8AzIEIQCUAH8AcgBcAC8AtgAYALoAuABBA00AcgAYAB8ATAFqAVUAmQCaAJoAmACyAAQAeABpABQAVwBuAM4AtAZUArgAZwUOAWUA5wAABMv+UgBa/6YAmf9nAG7/kgAt/9QAh/98ALgAqADlAI8AqAGF/nsAcAAeANkA3gFMBUYCzwVG/y0CigLZAlMClgC3AAAAAAAAAAAAAAAAAAABJQEYAOoA6gCuAAAAPgW7AIoE1wBTAD//jP/VABUAKAAiAJkAYgBKAOQAbQDuAOUASAPAADP+TgKx/0YDcAB5Bd8AUf+n/x8BCgBo/2wATwC8AKUHBQBhBysA7QSwAdIAtgB7AGUCUv90A2X+aQCUAI8AXABAAIYAdQCJAIlAQ1VUQUA/Pj08Ozo5ODc1NDMyMTAvLi0sKyopKCcmJSQjIiEgHx4dHBsaGRgXFhUUExIREA8ODQwLCgkIBwYFBAMCAQAsRSNGYCCwJmCwBCYjSEgtLEUjRiNhILAmYbAEJiNISC0sRSNGYLAgYSCwRmCwBCYjSEgtLEUjRiNhsCBgILAmYbAgYbAEJiNISC0sRSNGYLBAYSCwZmCwBCYjSEgtLEUjRiNhsEBgILAmYbBAYbAEJiNISC0sARAgPAA8LSwgRSMgsM1EIyC4AVpRWCMgsI1EI1kgsO1RWCMgsE1EI1kgsJBRWCMgsA1EI1khIS0sICBFGGhEILABYCBFsEZ2aIpFYEQtLAGxCwpDI0NlCi0sALEKC0MjQwstLACwFyNwsQEXPgGwFyNwsQIXRTqxAgAIDS0sRbAaI0RFsBkjRC0sIEWwAyVFYWSwUFFYRUQbISFZLSywAUNjI2KwACNCsA8rLSwgRbAAQ2BELSwBsAZDsAdDZQotLCBpsEBhsACLILEswIqMuBAAYmArDGQjZGFcWLADYVktLEWwESuwFyNEsBd65BgtLEWwESuwFyNELSywEkNYh0WwESuwFyNEsBd65BsDikUYaSCwFyNEioqHILCgUViwESuwFyNEsBd65BshsBd65FlZGC0sLSywAiVGYIpGsEBhjEgtLEtTIFxYsAKFWViwAYVZLSwgsAMlRbAZI0RFsBojREVlI0UgsAMlYGogsAkjQiNoimpgYSCwGoqwAFJ5IbIaGkC5/+AAGkUgilRYIyGwPxsjWWFEHLEUAIpSebMZQCAZRSCKVFgjIbA/GyNZYUQtLLEQEUMjQwstLLEOD0MjQwstLLEMDUMjQwstLLEMDUMjQ2ULLSyxDg9DI0NlCy0ssRARQyNDZQstLEtSWEVEGyEhWS0sASCwAyUjSbBAYLAgYyCwAFJYI7ACJTgjsAIlZTgAimM4GyEhISEhWQEtLEuwZFFYRWmwCUNgihA6GyEhIVktLAGwBSUQIyCK9QCwAWAj7ewtLAGwBSUQIyCK9QCwAWEj7ewtLAGwBiUQ9QDt7C0sILABYAEQIDwAPC0sILABYQEQIDwAPC0ssCsrsCoqLSwAsAdDsAZDCy0sPrAqKi0sNS0sdrgCIyNwECC4AiNFILAAUFiwAWFZOi8YLSwhIQxkI2SLuEAAYi0sIbCAUVgMZCNki7ggAGIbsgBALytZsAJgLSwhsMBRWAxkI2SLuBVVYhuyAIAvK1mwAmAtLAxkI2SLuEAAYmAjIS0stAABAAAAFbAIJrAIJrAIJrAIJg8QFhNFaDqwARYtLLQAAQAAABWwCCawCCawCCawCCYPEBYTRWhlOrABFi0sS1MjS1FaWCBFimBEGyEhWS0sS1RYIEWKYEQbISFZLSxLUyNLUVpYOBshIVktLEtUWDgbISFZLSywE0NYAxsCWS0ssBNDWAIbA1ktLEtUsBJDXFpYOBshIVktLLASQ1xYDLAEJbAEJQYMZCNkYWS4BwhRWLAEJbAEJQEgRrAQYEggRrAQYEhZCiEhGyEhWS0ssBJDXFgMsAQlsAQlBgxkI2RhZLgHCFFYsAQlsAQlASBGuP/wYEggRrj/8GBIWQohIRshIVktLEtTI0tRWliwOisbISFZLSxLUyNLUVpYsDsrGyEhWS0sS1MjS1FasBJDXFpYOBshIVktLAyKA0tUsAQmAktUWoqKCrASQ1xaWDgbISFZLSxLUliwBCWwBCVJsAQlsAQlSWEgsABUWCEgQ7AAVViwAyWwAyW4/8A4uP/AOFkbsEBUWCBDsABUWLACJbj/wDhZGyBDsABUWLADJbADJbj/wDi4/8A4G7ADJbj/wDhZWVlZISEhIS0sRiNGYIqKRiMgRopgimG4/4BiIyAQI4q5AsICwopwRWAgsABQWLABYbj/uosbsEaMWbAQYGgBOi0ssQIAQrEjAYhRsUABiFNaWLkQAAAgiFRYsgIBAkNgQlmxJAGIUVi5IAAAQIhUWLICAgJDYEKxJAGIVFiyAiACQ2BCAEsBS1JYsgIIAkNgQlkbuUAAAICIVFiyAgQCQ2BCWblAAACAY7gBAIhUWLICCAJDYEJZuUAAAQBjuAIAiFRYsgIQAkNgQlm5QAACAGO4BACIVFiyAkACQ2BCWVlZWVktLLACQ1RYS1MjS1FaWDgbISFZGyEhISFZLQAAAAIBAAAABQAFAAADAAcAACERIRElIREhAQAEAPwgA8D8QAUA+wAgBMAAAAUAd//KBp8F0wALABcAGwAnADMBB0AKkBmQGgJoCBobG7gCmkAPGBkUGBgZGBsVDxkaMSsSvAKfAAkBZQAMAp9ACwMaGRkDARsYGCUovAKfAB8BZQAuAp+yJQscvAKaACsBAAAxApqzIqw1BrwCmgAVAQAADwKaQAkgAAEAdTRXWhgrEPZd7fTtEPbt9O0AP+397RA8EDw/PBA8EO397QEREjk5ERI5OYcuK30QxDEwGEN5QFIBMykeKx8AMyAxHwEtJisfAC8kMR8BDQIPHwAXBBUfAREKDx8AEwgVHwEqHSgfATIhKB8BLCcuHwAwIy4fAA4BDB8BFgUMHwEQCxIfABQHEh8AACsrKysrKysrASsrKysrKysrgQFdEzQ2MzIWFRQGIyImASIGFRQWMzI2NTQmAwEzAQE0NjMyFhUUBiMiJgEiBhUUFjMyNjU0Jneeloq1t4aFsQE5Q1laQkRZWkIDIpL84QHlnpeKtbeHhbEBOkRZWkJFWVoEWp3cxb+6ycYBxXSbjXN0mo5z+nMGCfn3AY6e28W/usnHAcR0m4x0dJqOcwABAHz+UQJgBdMAEAA9QAonDwEAEBIHCBAQuAEzswCfDgi4ATNAEQefDl4AAxADIAMDA6wRnYwYKxD2Xf327RD27QA/PD88MTABXQEmAhE0NzY3MwYHBgcGFRABAd+Vzk1avIF5Jz0jKwEr/lG8AfgBDu7a/fvQWYqWu73+H/4gAAEAfP5RAmAF0wAQAGVADCgCKBACCQoQAQASCbgBM7MKnwMBuAEztACfA14OuP/wtBAQAlUOuP/4tA8PAlUOuP/ktA0NAlUOuP/sQA8KCgJVDw4fDgIOrBKdjBgrEPZdKysrK/327RD27QA/PD88MTABXRMjABE0JyYnJiczFhcWFRAC/YEBKysiPSd6gbxaTc/+UQHgAeG8uZaKWtL7/dru/vL+CAABAHIA7QQ6BLYACwA4QB8AbgkC+QgDbgUHBgluCgQK+QUBbj8CTwICAhkMV1oYK04Q9F1N9DztPBDkPDwAL/Q8/Tz0MTAlESE1IREzESEVIRECAf5xAY+qAY/+ce0BkqgBj/5xqP5uAAEAqv7eAYMAzQAKAE61CgMAB6sGuAFQQCYBAzwCAgEKATwACgIDAQM8AAY4BzpPAF8AbwB/AKAABQCgC6GYGCsQ9F305BDtPBA8AD/tPBA8EO0Q/e0BERI5MTAzNTMVFAYHJzY2N7bNUFcyOTYDzc1xiyZNGWFbAAEAQQG4AmoCbQADACxAGXACcAMCTQFNAgIBIwACGgVwAAEAGQRwjRgrThDkXRDmAC9N7TEwAHEBXRM1IRVBAikBuLW1AAABALoAAAGHAM0AAwAlQBgCPAAKAjxfAG8AfwCvAASgAAEAoAShmBgrEPZdXe0AP+0xMDM1MxW6zc3NAAABAAD/5wI5BdMAAwBTuQAD/96yFDkCuP/eQCAUOZcDAQIDnwOvAwIDdgABFAAAAQIBAAMACgPoAALoAbgBqbUAAASzehgrEDwQ9O0Q7QA/PD88hwUuK119EMQxMAFdKysVATMBAamQ/lgZBez6FAAAAgBV/+cEEQXAABAAHQFVsQICQ1RYQAoaHgQFFB4NDRcJuP/otA8PAlUJuP/oQBkNDQJVCREADA8PAlUAFgwMAlUADA0NAlUALysrK80vKyvNAD/tP+0xMBuxBgJDVFhAChoeBAUUHg0NFwm4//S0Dw8GVQm4/+a0DQ0GVQm4/+5AGQsLBlUJEQAQDQ0GVQAQDAwGVQAQCwsGVQAvKysrzS8rKyvNAD/tP+0xMBu0BiAZEBy4//CyAiALvv/gABb/4AAS/+AAD//gQGIEBocCiAuID8kOBQkHCxgCRRNMFUoZQxtUE1wVXBlSG2sHawtjE2wVaxlgG3kCdwZ2C3oPhwaYB5YQyRjaAtYG1gvbDxoaHgQFFB4NDRdzCUAhIzQwCQEACRAJAgmQHxFzALj/wEAOISM0IABAAAIAkB7HixgrEPZdK+0Q9l1xK+0AP+0/7TEwAV1xAF0AODg4ODgBODg4WVkTEBI2MzIWFhIVEAIGIyInJhMQFjMyNhEQJiMiBwZVa9OgdrJ0QmrTodR5kbmpfHypqX58Sl0C0wEEAT2sX7P+/9r+/v7DrZi3AZ3+l+/wAWgBau5phgAAAQDfAAAC+wXAAAoAr0AgA0ANETRrBH8CjwKZCASsBAEJAAYFAgMJBQEMAgHKCgC4/8BACiEjNDAAASAAAQC4/+C0EBACVQC4/+pAEQ8PAlUAHAwMAlUADg0NAlUAuP/wQBkPDwZVABAMDAZVABANDQZVABoMBUANDzQFuP/AQA4hIzQwBQEgBUAFAgUZC7oBPAGFABgrThDkXXErKxD2KysrKysrK11xKzxN/TwAPz8XOQEROTEwAV0AXSshIxEGBgc1NjY3MwL7tEHTVJfiL3QEez58H65Hyl8AAAEAPAAABAcFwAAeAcexBgJDVFhACREQDRgTEwZVDbj/9LQREQZVDbj/7kAJEBAGVQ0eFAUeuP/oQBcTEwZVHh4REQZVHhwOEAZVHgwNDQZVHrgCu0AMAgoXFyAfEBECAiAfERI5L9TNERI5L80AL+0rKysrP+0rKyvEMjEwG7ECAkNUWEAJERANDBISAlUNuP/0QAkPEQJVDR4UBR64/+BACxITAlUeFA8RAlUeuAK7sgIKF7j/6LQLCwJVF7j/7EAODQ0CVRcXIB8QEQICIB8REjkv1M0REjkvKyvNAC/tKys/7SsrxDIxMBtANjsFOwa7Bb8GuwfHCMkcB0kMWQxUDmsMZA56EnoTiRK8EuUa5RvwGgy/C7cTAhsQHBAdEB4QBr7/8AAH/+AACP/wAAn/8EAaHgoQCAYGyhwaFBwcGggcGgMBAggaHAMNHhC4AqSzTxEBEbgBGLUNHhQFAB64ArtADwECDApzF9MAAAFAISM0AbsCgQAgABABOEAMEbU/Al8CbwJ/AgQCugIkAB8Bj7GLGCsQ9l307RD2KzwQ9O0APzz9PD/t/V3kERIXOQEREhc5hw4uKw59EMQBERI5MTAAODg4OAE4ODg4AF0BXXJZWSUVISY3NjY3NjY1NCYjIgYHJzY2MzIWFRQGBgcGBgcEB/w3Ahclo5rvqJl7gpwBuRP40dP2SKfColwera1BPGPAfsTlZmuTnIoTz9nqrViqvKSIYTEAAQBW/+YEFgXAACsBWbECAkNUWEALGRhADQ0CVRgcAAG4/8BAKwwNAlUBKSMKDQ8MDx4KCikVHhwEHikcBSkNIw0MGBkBABIgEAwMAlUgBya4/+i0DA0CVSYvK80vK80vzS/NLwASOT8/EO0Q7RI5L+3GEMYSORDEKzIQxCsyMTAbQCgFDRYNRQ2GDQRFEVcRdhsDUhZsEGoUZBZ1DXkUhg2KFIkbpQ0KBSADuP/gQAsLDA0OBAcBIw0MAbgCpLNAAAEAuwEYACkADQE1tAwMFQQYugKkABkCaEAnFR4cBQQeKQ0Sc18gbyACIBgNDQZVIIAHcyZAISM0MCYBACYQJgImuP/0tw0NBlUmkC0YuAE4shnTAboBOAAA/8BACyEjNCAAQAACAJAsuAGSsYsYKxD2XSvt9O0Q9itdcSvt9Ctd7QA/7T/t/eQREjkv7RD9XeQREjkBERIXOTEwATg4AV0AXQFxWRM3FhYzMjY1NCYjIgc3FjMyNjU0JiMiBgcnNjYzMhYWFRQGBxYWFRQAIyImVrQflWt/r6J9M0wUEgtzuIZqaYwUtCHqrnjKa2ZkgpD+6NbB/wGDGJmHsIJ8oRSeAnh9Y4KEhCC1x2eyZF+cLh69jsD+9eYAAgAaAAAEEAW6AAoADQEmQDYSWAxoDJoMqQzJDAVMA0wNlAQDEgECCAAMBgMHBQoLAwcADAwNDcoDBBQDAwQDDQACDA0EBwO7ArsACAACAaBACgAEBAAMDADKCgS4Ama3BQUKQB0fNAq4/+C0EBACVQq4/+a0DQ0CVQq4/+60DQ0GVQq4ATdADQdAIiM0B4AhNQeQDwK4/8BACw0UNAACEAIgAgMCuP/gtA0NAlUCuP/ktg0NBlUCtQ64AYyxixgrEOwrK10rEPYrK/QrKysrPBDmEP08AD8/EPQ89jwROTkBERI5OYcuKwR9EMQPDw8xMAFDXFi5AA3/3rISOQ24/9RACzM5AyItOQMEHR08KysrK1ldAF1DXFhAFAxACzkMgFA5DEAmOQwiHDkMQC05KysrKytZIREhNQEzETMVIxEDEQEClv2EAp2Txsa0/jUBX6UDtvxKpf6hAgQClf1rAAEAVf/nBCEFpgAeAVaxAgJDVFi5AAH/wEANDQ0CVQEcDgoeFRUcErgCu0ALDwQEHhwNDgEABxi4/+q0Dw8CVRi4/+q0DQ0CVRgvKyvNL80vAD/tP+0SOS/9xBDEKzEwG0ApEgwNDQZVDwwNDQZVSxp5HYodlhOnE8MM1gzbGwgJExgOKhoDCTAFMAu6/+AAA//gQBATChUSExPKDg8UDhMUDg8NuAKkQBMOCh4VQA6gDgIODg9AFQEVFRwSuAK7tw8EAdNAAAEAuAEYQCAEHhwNEV8QbxB/EI8QBBCAB3MYQCEjNDAYAQAYEBgCGLj/9LcNDQZVGJAgErwBNQAPAZUADQE4sg61AboBOAAA/8BACyEjNCAAQAACAJAfuAGSsYsYKxD2XSvt9O307RD2K11xK+30XTwAP+39XeQ/7RI5L10ROS9dEO0Q5IcILisFfRDEABESOTEwATg4ODgBcV0rK1kTNxYWMzI2NTQmIyIGBycTIRUhAzYzMgAVFAcGIyImVb0VmWyCtK2MV4woqY4C2f23T4SRwAEIdI30yP0BgBCKi8SimrJPPxYC8az+dlz+9tHHkbLgAAACAE3/5wQVBcAAHQAqAU+xAgJDVFhAHw8BHwFfAQMBGygeQA0BDQ0UBR4bBSIeFA0KHgEAJRC4//RAGQ0NAlUQHhcQDw8CVRcQDAwCVRcMDQ0CVRcvKysrzS8rzdTNEMUAP+0/7RI5L13tEMRdMTAbQC1rGQFEB0AVRBlEIFoSVCBrA2QHZAhqEmQgdAh1HIUIhhzWCNQWEQcgDQ0GVSe4/+C0DQ0GVSO4/+BACw0NBlUhIA0NBlUHuP/gtCcgIyAhuP/gQBEoHkANUA0CDQ0UGwHTXwABALgCaEAJBR4bBSIeFA0BuAE4QBIAtSVzEEAhIzQwEAEAEBAQAhC4//C3DAwGVRCQLAq6ATgAHgE5QBY/F18Xbxd/FwQXFgwMBlUXFg0NBlUXuAIksyvHixgrEPYrK13t7RD2K11xK+307QA/7T/t/V3kERI5L13tMTABODg4OCsrKysBXQBdWQEHJicmIyIHBgYHNjYzMhIVFAYGIyIAERA3NjMyFgEUFhYzMjY1NCYjIgYD+7MYLElrVkFVYgJBvGe0/XfQhOH+5J2J6K3d/TdPjk5ypKJ7eqoEUw5qME0wPu7cY2D+99KK7X4BSwF8AanBqML83V2qWbiemK+vAAEAYQAABBYFpwANAHBADsQNAQQNAQQCCAQJAw0AuAK7QDACAQQJDA1zAwMCQCEjNE8CXwJvAgMCGg8IcwnrAE8BXwFfAgM/AV8BbwF/AQQBGQ64AZKxixgrThD0XXE8TfTtThD2cSs8TRDtAD8/PP08ORE5ARESOTEwAXFdEzUhFQYAAwYHIzYSEjdhA7WM/u1LNg+5A4LziQT6rYyV/hL++7jbrQHqAcecAAADAFP/5wQZBcAAFwAjADACALECAkNUWLQMABseLrj/wEAXExMCVS4uEiEeBgUoHhINHgkMDAwCVQm4//S2DQ0CVQkrD7j/8LQPDwJVD7j/6LQLCwJVD7j/6LYNDQJVDxgDuP/wtBAQAlUDuP/wtA8PAlUDuP/0QBkNDQJVAyQVDAsLAlUVDAwMAlUVDA0NAlUVLysrK80vKysrzS8rKyvNLysrzQA/7T/tEjkvK+05OTEwG7EGAkNUWLceCQwMDAZVCbj/9LYNDQZVCSsPuP/ktA8PBlUPuP/ktg0NBlUPGAO4//C0Dw8GVQO4//xAIg0NBlUDJBUMDAwGVRUMDQ0GVRUMABseLi4SIR4GBSgeEg0AP+0/7RI5L+05OQEvKyvNLysrzS8rK80vKyvNMTAbQDc1FgEpFkkWSSbmDOkwBQkwAX0AfQF8BHQIcQtyDHUNeheLAIoBjASGCIELhAyGDY0XzBHGExIiuP/gshwgGrj/4LIgIC+4/+CyLSAmuP/gQB4pIAwAHhgADBseLqAuAS4SIR4GBSgeEg0ec78JAQm4AmdAECtzD0AgIzQwDwEADxAPAg+4AZG2MhhzsAMBA7gCZ7IkcxW4/8BADiEjNCAVQBUCFZAxx4sYKxD2XSvt9F3tEPRdcSvt9F3tAD/tP+0SOV0v7Tk5ARESOTkxMAE4ODg4ODg4OAFdcnEAcVlZASYmNTQ2MzIWFRQGBxYWFRQAIyIANTQ2ExQWMzI2NTQmIyIGAxQWFjMyNjU0JiMiBgFqcGzmv8Dqa22Hjf722dn+9pFihmtohYlmZ4g6SZBTgaitgn+nAxspmGqg2t+gZpcpLMSIvP8AAQHAj8EBVGiEg19jh4T8/02QT6aAgqqoAAACAFX/5wQZBcAAHgAqAa6xBgJDVFi3Cx8YAQAlERi4//a0Dw8GVRi4//S0DQ0GVRi4//BAKAwMBlUYEQwNDQZVERAMDAZVERgRLCsLKB4PDh8OTw4DDg4UAFABAQG4/8BADRARBlUBBB4cDSIeFAUAP+0/7cQrXTISOS9d7TIBERI5OS8rKy8rKysQzdTNEN3FMTAbsQICQ1RYtwsfGAEAJREYuP/qtA8PAlUYuP/qQCoNDQJVGBEMDAwCVREYESwrCygeDw4fDk8OAw4OFABQAQEBBB4cDSIeFAUAP+0/7cRdMhI5L13tMgEREjk5LysvKysQzdTNEN3FMTAbQDQ6GkwWQCNbFlcjZgNsFm0aZyN6Gn0ejBqLHpoWqRq8GuoW5iD2IBM9Fp4WrRYDOilkBgInuv/gACP/4EAYISAGICgeTw5fDgIODhwiHhQFAdNQAAEAuAJotAQeHA0fugE5AAsBOEARGEAhIzQwGAEAGBAYAhiQLAG4ATi0ALUlcxG4/8BADiEjNCARQBECEZArx4sYKxD2XSvt9O0Q9l1xK+3tAD/t/V3kP+0SOS9d7TEwATg4ODgAXXEBXVlZEzcWFjMyPgI1NCcGBiMiAjU0ADMyFhIREAIGIyImATQmIyIGFRQWMzI2cK0WfGFTfVA2ATa7bbb8AQfGj+17evGirNoCy6V0eLKpfH2hAVMQem5Mf9hwDBhWawEI2N8BEJr+4/7y/uf+s66/AzSbtsScjK+vAAACALkAAAGGBCYAAwAHADhAIAQFAAYHCQIGPAQDPAEGBAoCPC8APwACIAABAKEIoZgYKxD0XXHtAD8/7RDtARESOTkSOTkxMBM1MxUDNTMVuc3NzQNZzc38p83NAAIAcgGhBDoEBgADAAcAR0AnBQYBBAcJACUDASUDAgclBAQGJTACAZ8CzwICAr8FABoJARkIV1oYK04Q5BDmAC9N7V1x7TwQ7RA87RDtARE5ORE5OTEwASE1IREhNSEEOvw4A8j8OAPIA16o/ZuoAAACAFoAAAQMBdMAHgAiAIRAL4waixsCfBp8GwJiGmUbAmsMYQ4CWgxUDgI2DkQOAhsZCAcEABAnEREADSkUAR4AuAKvQCMhIiE8HwofPCIiIDwhIR4AXh5uCl4XaiQQXiARARFqI1daGCsQ9l3tEPbt9O0QPBDtPBD9AD/tPBD2PD/tEjkv5BEXOTEwAV1dXV0AXV0BJjU0NzY3PgI1NCYjIgYHJzY2MzIEFRQGBw4CBwM1MxUB2AEeFjEkuzikd3OaGLkZ98vXAQBag1g2GgK4zQFpJBJqTTo7K6ViOmmfkJkWzdrqpmCidE5KYGz+l83NAAL//QAABVkFugAHAA4BZ7YBDg8QAlUCuP/ytA8QAlUCuP/4tA0NBlUCuP/0QFkMDAZVCQwMDAZVBQwMDAZVLxAwEGcIaAlgEIgDkBDJBcYGwBDwEAsIBVkBVgJQEGgLsBDzDPMN8w4JBAwEDQQOAwsKCQUEBAwNDggGBwcMCQUECAYMBwEAALj/+EAPDAwCVQAgBwwUBwcMAgMDuP/4QBUMDAJVAyAEDBQEBAwJHgUFCB4GAwa4AnBACQAIDOlAAgECAroBCwABAQtAEgwgAGUHA1JQBM8E3wQDkAQBBLgBAUALUAzAB98MA5AMAQy4AQFAEA8HzwcCfweABwIHkw/W1xgrEPRdcRn0XXH0XXEY7RDtGhkQ7e0AGD88Gu0/5DwQ7TwQ7YcFLisrfRDEhy4YKyt9EMQBERI5ORE5OYcQxMQOxMSHBRDExA7ExDEwAUuwC1NLsB5RWli0BA8DCAe6//AAAP/4ODg4OFkBcnFdKysrKysrIwEzASMDIQMTIQMmJwYHAwIz0QJY3av9m6HZAfGZRiIcMwW6+kYBvP5EAloBlrl3jYsAAAMAlgAABOkFugARAB0AKgETuQAE//RARwsLBlUEBEYjViNmI3MJhAkGaRp1BXAJcwuDBYMLBicWCQMYJyoeFh0JCRMSHioqKSkAHB0eAgECHx4eEQAIGCYGDBAQAlUGuP/mQDMPDwJVBhINDQJVBgYMDAJVBggLCwZVBgwMDAZVBhQNDQZVBlQlJgwcEBACVQwKDQ0CVQy4//RAFQsLBlUMGiwdHiABIAABACAQEAJVALj/9rQPDwJVALj/9rQNDQJVALj/+rQMDAJVALj/+rQMDAZVALj/8EAKDQ0GVQBdKztcGCsQ9isrKysrK108/TxOEPYrKytN7fQrKysrKysr7QA/PP08Pzz9PBI5LzwQ/Tw5LxE5ERI5ARIXOTEwAV0AXSszESEyFhYVFAYHFhYVFA4CIwEhMjc2NjU0JiYjIREhMjc+AjU0JiYjIZYCJqjLc2ZnhY9XgMGM/pMBPYE4SktGgp7+2wFtXiZDWjpUlYz+rQW6WbllXqYzJ7yAZ7FgMQNSERZmTUlvKfugBww4a0ZSeTEAAAEAZv/nBXYF0wAdANO1YwJqHQIBuP/otAsLBlUAuP/oQF8LCwZVIAAyDWMAcAB0HYAAhB2QAJoFqwOlDbkDtA3HDdAA5B3zHREOEh0RHR0DKgYoESocIB9HDVYUVxVWGWgFax17EosSmgOZDpocqAGkAqgR1Q4TABQAGhAUEBoEArj/3rIoOQG4/8BALSg5EA8AAQQbEx4MAxseBAkQJg9KACYgAQEBGh8XJiAIAQgMCwsGVQgZHmNcGCtOEPQrXU3tThD2XU3t9O0AP+0/7REXOTEwASsrXV1xAF0rKwFyARcGBCMiJAI1NBIkMzIEFwcmJiMiBgIVFBIWMzI2BLTCPf7D5e3+15uvAUPC3AEsO78zwpOp41xt5oaj4gICMe/7wQFu0uUBVbHgyy2gkqL+75G7/umKvAAAAgCeAAAFWgW6AA8AHQDlQC8gHwFDCBwdHgIBAhEQHg8ACBcmIAkBH0ANDQJVCSAQEAJVCQoPDwJVCRgNDQJVCbj/9EAVDAwGVQkaHx0QIAEgAAEAIBAQAlUAuP/2tA8PAlUAuP/2tA0NAlUAuP/6tAwMAlUAuP/3tAwMBlUAuP/4QAoNDQZVAF0eO1wYKxD2KysrKysrXTz9PBD2KysrKytd7QA/PP08Pzz9PDEwQ3lANgMbBwgGCAUIBAgEBhkYGhgCBgsKDAoNCgMGFRYUFhMWAwYbAxchARIOFyEBGAgcIQEWChEhACsrASsrKioqKoEBXTMRITIXFhcWEhUUAg4CIyUhMjY3NjY1NCYnJiMhngH5q1p+WXRzTnqRzYX+sQE5kaUxRU2XbE6t/swFuhUdTGL+z8Sn/v6pYTKtNjFF6abm9yoeAAEAogAABOgFugALAJVAFQYFHggIBwcAAwQeAgECCgkeCwAIB7j/wEAdEBI0B1QDSiAKIA0CChoNBAkgASAAAQAgEBACVQC4//a0Dw8CVQC4//a0DQ0CVQC4//q0DAwCVQC4//q0DAwGVQC4//BACg0NBlUAXQw7WxgrThD0KysrKysrXTxN/TxOEPZdTfTkKwA/PP08Pzz9PBI5LzwQ/TwxMDMRIRUhESEVIREhFaIEJPyeAyv81QOEBbqt/j+s/g2tAAABAKgAAASFBboACQCNQCsGBR4ICI8HAQcHAAMEHgIBAgAIB5wgAiALAgIaCwQJIAEgAAEAIBAQAlUAuP/2tA8PAlUAuP/2tA0NAlUAuP/6QAsMDAJVAAwLCwZVALj//rQMDAZVALj/8EAKDQ0GVQBdCjtcGCtOEPQrKysrKysrXTxN/TxOEPZdTeQAPz88/TwSOS9dPBD9PDEwMxEhFSERIRUhEagD3fzlArD9UAW6rf46rf1mAAEAbf/nBbkF0wAlARNAGhsUGxUCYCcBXggTARIDJCQAIRIXAiUAHgIBuP/AQCAMDAZVAQEGFx4OAyEeBgkBASYnJSQgAwMgAiAnYAIDArj/5LQPDwJVArj/8rQNDQJVArj/2rQMDAJVArj/9EAbDAwGVQJygCcBJx0mIAoBChAMDAZVChkmY1sYK04Q9CtdTe1NEF32KysrK108TRD9PBESOS8AP+0/7RI5Lys8/TwREjkREjkBERI5EjkxMEN5QEQEIxscGhwZHAMGDCYQJRUmHyYIJQQmIyUYDR0hABYPEyEBERIUEyAHHSEAIgUlIQEcCxchARQRFyEBHgkhIQAkAyEhAAArKysrASsrEDwQPCsrKysrKysrKyqBAV0AXQE1JREGBCMiJAI1NBIkMzIEFhcHLgIjIgYGBwYVFBIEMzI2NxEDTAJtj/7QoNj+n7SzAVDbnwEBkiavIWK2b4XCdyE4hwECkX7wPgI/rAH94HJzuQFe2NYBc7RnuJQwcIBNUYRPiJ/E/viAYTcBEQABAKQAAAUiBboACwDYuQAN/8BAGhMVNAQDHgkKoArQCgIKBQICCwgIBQggBwcGuP/utA8PAlUGuP/yQAsNDQJVBhAMDAJVBrj/4EAYCwsGVQYBDAwGVQZdgA0BDQILIAEgAAEAuP/AQAoTFTQAIBAQAlUAuP/2tA8PAlUAuP/2tA0NAlUAuP/6QAsMDAJVAAgLCwZVALj/97QMDAZVALj/+EAWDQ0GVQBdDCANASANUA1gDXANBDtZGCtdcRD2KysrKysrKytdPP08EF32KysrKys8EP08AD88Pzw5XS88/TwxMAErMxEzESERMxEjESERpMIC+sLC/QYFuv2mAlr6RgKz/U0AAQC/AAABgQW6AAMAzLUBAgAIAgW4/8CzOD00Bbj/wLMzNDQFuP/Asy0wNAW4/8CzKCk0Bbj/wLMjJTQFuP/Asx0eNAW4/8CzGBo0Bbj/wEAqDRA0IAWQBa8FAwMgAQAAjwCgALAABC8AQABQAN8A8AAFEiAAjwCQAAMFuP/AQAsNDQJVABgQEAJVALj/7LQPDwJVALj/7rQNDQJVALj/9kAQDAwCVQAgCwsGVQCiBNZZGCsQ9isrKysrK11DXFiygAABAV1ZcXI8/V0rKysrKysrKzwAPz8xMDMRMxG/wgW6+kYAAQCWAAAEKgW6AAUAbUAMAQIEAx4FAAggBAEEuAKnQA8HAgMgASAAAQAgEBACVQC4//a0Dw8CVQC4//a0DQ0CVQC4//q0DAwCVQC4//a0DAwGVQC4//hACg0NBlUAXQY7XBgrEPYrKysrKytdPP08EOZdAD88/Tw/MTAzETMRIRWWwgLSBbr6860AAQCYAAAGDwW6ABAC5LECAkNUWLkACP/2QAsMDAJVCA4NEQJVArj/7rQNEQJVBbj/7kAoDRECVQwSDAwCVQUPDAMJAAECCAkLDgAICQIKCwYQEAJVCxANDQJVC7j/+rYMDAJVCxAAuP/mtBAQAlUAuP/4tA8PAlUAuP/8tA0NAlUALysrK80vKysrzQA/P8DAENDQwBESFzkrKzEwASsrKwAbsQYCQ1RYQB8HIAsLBlUGIAsLBlUDIAsLBlUEIAsLBlUFIAsLBlUIuP/yQCMLCwZVAgwLCwZVAwYMDAZVAg4MDAZVCQwMDAZVCgwMDAZVB7j/+LQNDQZVCLj/+EAfDQ0GVSYFAQwgChI0DyAKEjQPBQwDAAEOCwAICAECCrj/7rQLCwZVCrj/7rQMDAZVCrsCVgASABACVkANAAwLCwZVAAYMDAZVALj/+LQNDQZVAAEvKysr9C/0KysAPzw/PDwREhc5KytdMTABKysrKysrKysAKysrKysbQH8AAg8IFAIbCAR2DIYMyAwDCQxJDEkPAykEJQ0sDlgDWwR2DXgOhw0ICwIFCDkNNg5PAksDRAdACE0NQg4KmAKZA5YHlgioA6cHBhICDw4OMAUCFAUFAggMDQ0wBQgUBQUIDFIPUgFAAQICCAgJCgsLDQ0ODhAACAkCYBKAEgISugKoAA0BMbIFIAi4ATFACgwJCiBADH8LAQu6AlYADgELsgUgArgBC0AJDwEAIA9wEAEQuAJWtyAFYAWABQMFuAKosxE7WRgrGRD0XfRdPBj9PBDtGhkQ7fRdPBoY/TwQ7RoZEO3kXQAYPz88PBA8EDwQPBA8EDwQPBoQ7e2HBS4rh33Ehy4YK4d9xDEwAEuwC1NLsB5RWli9AAz/+wAI/9YAAv/WODg4WQFLsAxTS7AoUVpYuQAN//ixDgo4OFkBQ1xYuQAN/9S2ITkOLCE5Dbj/1LY3OQ4yNzkNuP/UtS05DiwtOSsrKysrK1lycV0AcV0BXVlZMxEhARYXNjcBIREjEQEjARGYASQBWzAWGTUBXwEFu/5Wr/5YBbr78pFIUJsD/PpGBMv7NQTg+yAAAQCcAAAFHwW6AAkBfbESC7j/wEAKExU0CBgMFgJVA7j/6EAhDBYCVQgCAwMgBwgUBwcIAgcDAwgJBAICCQcIBAMgBgYFuP/stA8PAlUFuP/yQAsNDQJVBRIMDAJVBbj/90AaCwsGVQVdIAsBIAtQC2ALcAuACwULCAkgAQC4/8BADRMVNCAAAQAgEBACVQC4//a0Dw8CVQC4//a0DQ0CVQC4//pACwwMAlUABAsLBlUAuP/3tAwMBlUAuP/4QAoNDQZVAF0KO1kYKxD2KysrKysrK10rPP08EF1x9CsrKys8EP08AD88PzwSOTkBETk5hwQuK4d9xLEGAkNUWLkAA//gtwwRNAggDBE0ACsrWTEwKysBK0NcWLQIQEY5A7j/wLZGOQhAMjkDuP/AtjI5ByIZOQK4/962GTkHIjI5Arj/3rYyOQciIzkCuP/eQAsjOQcOFDkHDhM5Arj/9LYTOQcOHTkCuP/0th05Bw4VOQK4//ixFTkrKysrKysrASsrKysrKwArKysrWTMRMwERMxEjARGcxwMCusf8/gW6+4EEf/pGBID7gAAAAgBj/+cF3QXUAA4AGwDKQFAaDwEUEBQUGxcbGwQEEAQUCxcLGwSpF7YOxg4DFxcYGwIgHUARTxNPF0AaWAVYCVcQVRFfE1oXXxhWGlcbixeZAhAZHgMDEh4LCRUmIAcBB7j/6LQQEAJVB7j/7rQNDQJVB7j/8LQMDAJVB7j/6rQLCwZVB7j/9LQNDQZVB7j/+kAhDAwGVQcagB0BHQ8mIAABAAYLCwZVAAYMDAZVABkcY1wYK04Q9CsrXU3tThBd9isrKysrK11N7QA/7T/tMTABXXEAXV1dcRMQACEyBBIVFAIEIyIkAjcQADMyABE0AiYjIgBjAYgBNssBRqu0/ra/z/66qMgBHdfbARt56ZHO/tcCygFtAZ3C/qXc3/6gtcgBWr7+9/7PATQBG7MBC5P+5QACAJ4AAAT9BboADQAYALJALGURaxQCSxBLFFsQWxQECwweDw4OABcYHgIBAgAIEiYICg0NAlUIEAsLBlUIuP/0QBsMDAZVCBogGgEgGgEaGA0gASAAAQAgEBACVQC4//a0Dw8CVQC4//a0DQ0CVQC4//pACwwMAlUADAsLBlUAuP/6tAwMBlUAuP/wQAoNDQZVAF0ZO1wYKxD2KysrKysrK108/TxOEHFd9isrK03tAD8/PP08EjkvPP08MTABXQBdMxEhMhceAhUUAiEhEREhMjY1NCYnJiMhngIpkk1sklnu/sn+iAF7vJ5dTDGE/okFug4SZbZtu/79/awDAYx/XIMVDQAAAgBY/44F7gXUABUAKAFoQJVfJp8mAhkYNxUCCxwEHwQjGxwUHxQjBioFLRcrJjsFPBc6JkwFTBdJJl0FVSNYJm8FewN6BYwDjAWVAJoDpACrA9UA1RblAOUX5RgaHAUrACoFOwUEXQWSGJYm1SYEJRYqJjQWOSZJGEkcRR9FI0smVghYEVUVWhxaHVYfVyBXImkFZhVrJnsmjhyOJtsY3CYZCxgBFbj/1LIbOQC4/9RAOBs5BBgUGCoFOgUEAgMWKAMHKCYYFgUABiEDExoFAigmGBYABSQeHg8DAggkHgcJGiYTGA8PAlUTuP/utA0NAlUTuP/otAwMAlUTuP/wtAsLBlUTuP/0tA0NBlUTuP/0QCUMDAZVE0oCGiAqgCoCKiEmIAsBCxgLCwZVCwYMDAZVCxkpY1wYK04Q9CsrXU3tThBd9k30KysrKysr7QA/7T8/7REXORI5ARESORIXOQARMxDJEMldMTABKytdXQBycV0BXXFyJRYXByYnBiMiJAI1NBIkMzIEEhUUAiUWFzYRNAImIyIAERAAMzI3JicE9YdyOZ6do8XH/ryvsAFFycsBRqtu/eaobat56ZHZ/uIBG9xoXFtlnV0rhzl7W8ABXNrZAWS6wf6l2rX+340vXZwBObIBCpP+1/7Z/uL+zic7GQACAKEAAAWtBboAGAAiAfxAIRILDgESNhxaH2YIbR8ECRANDQZVCBANDQZVBxANDQZVJLj/wLQMDAJVDbj/9LQMDAJVDLj/9LQMDAJVC7j/9LQMDAJVErj/4rMSGjQSuP/wsyInNBG4/+KzHSc0ELj/4rMdJzQPuP/isx0nNBK4/9izHSY0Ebj/4rMSGjQQuP/isxIaNA+4/+JASRIaNCUOShxKIFMLXBxtHHIJeA55D4UKiA+XDakPuA/oDucPEA4MDCARDxQREQ8RDwwJEhsCIRoWCgYSERANDAUYCQkWFxoZHhe4/8BAGQsLBlUXFwAhIh4CAQIAGBgPDw4IHiYOnAa4/+i0Dw8CVQa4//a0DQ0CVQa4/+BAIgwMAlUGBg0NBlUGXSAkcCSAJAMkIhggASAAAQAgEBACVQC4//a0Dw8CVQC4//a0DQ0CVQC4//pACwwMAlUABgsLBlUAuP/3tAwMBlUAuP/4QAoNDQZVAF0jO6gYK04Q9CsrKysrKytdPE39PBBd9isrKysZ5BjtAD88EDwQPD88/TwSOS8r/TwQPDkvEhc5AREXOYcOLisFfRDEMTABXSsrKysrKysrKysrKysAKysrXUNcWEAKCEAPOQ8QOhESOisrK1kBcUNcWLkADv/eQBoZOREiGTkSIhk5DkAcORAiFDkQIh85ECIVOSsrKysrKytZMxEhMhYWFRQGBxYXFhcTIwMuAicmIyMRESEyNjY1NCYjIaECisTMesrTTShVTP/0wlVuVy0hS+EBoYWWTpej/jAFuk/IeZzWHSUkTnX+cQExhIw4Cwf9dQMzN3lHaIYAAAEAXP/nBOsF0wAwAhVAJ2MDYwRzA3QEBCUnNQM5HEMDSQdMHUUfRCRGJ1MDWQdcHVcoiRMOI7j/8rQQEAJVJLj/8rQQEAJVJbj/8rQQEAJVJrj/8rQQEAJVJ7j/8rQQEAJVI7j/9rQNEAJVJLj/9rQNEAJVJbj/9rQNEAJVJrj/9rQNEAJVJ7j/9kBGDRACVSgNJiQCJAMnJTYPNCNEJUUvWiBWI1UlbAtqDWsOZhRlGHkLeg16D30QdSRzJYYDiguJDYoPjRCFJIMlkg2WD5YVHrEGAkNUWEAtISYSGyYaCSYpASYAACkaEgQyMSYAZQACAA0teRuJGwIbJRYNLR4nJQElBRYFuP/0QAwMDAZVBR4tCR4eFgMAP+0/7SsREjldERI5ERI5XRESOV0BERIXOS/tL+0v7S/tG0AtJSQODQsFIRwdHhsIBwYEAwIGASUkIg4NCwYFHhstGkAMDAJVjxoBGu0WAC0BuP/AQBIMDAJVEAEgAVABYAFwAZABBgG4AbBAEy0eHhYDBR4tCRsmGkoJJgApASm4/+q0Dg4CVSm4//RADQwMAlUpGjIhJhIBJhK4/+y0Dg4CVRK4//a0DQ0CVRK4//hADwwMAlUSVCAAAQAZMWNbGCtOEPRdTeQrKyvtEO1OEPYrK11N7fTtAD/tP+0Q/V0r5BD9XSv0ERIXOREXORESOTkBEhc5WTEwAF1xKysrKysrKysrKwFdcRM3HgIzMjY2NTQmJyYkJyYmNTQ2NjMyFhYXByYmIyIGFRQXFgQXFhYVFAYGIyIkJly3DV/IfW+qU1BcO/5sUWlnfvKUo/mGBboPramwoTk4AdlYgHqG+53H/vOZAdcQbo1XQnNERWcjF2ErN6Nlb8FkacyBDouOgVtPMzNrKDu1dnXPc3TpAAABADAAAAS6BboABwCJQA0FAh4EAwIACAcGBQQJuAJzsyAEAQS4AQG3BiABAi8DAQO4AQG1AQEgAAEAuP/oQAsQEAJVAAgPDwJVALj/8rQMDAJVALj/4rQNDQJVALj//LQMDAZVALj//rQNDQZVALgCc7MItpkYKxD2KysrKysrXTwQ9F08EP3kXeYQPBA8AD8/PP08MTAhESE1IRUhEQIT/h0Eiv4bBQ2trfrzAAABAKH/5wUiBboAFADZQAomD1gEWAjJCAQWuP/AQBYTFTQ0BDsIRgRKCHYPpgXoDwcMAAIRuAK7tAYJFCYCuP/stA8PAlUCuP/yQAsNDQJVAhAMDAJVArj/4EAcCwsGVQJdIBYBIBZQFgJgFnAWgBYDFg0mIAoBCrj/wEAKExU0CiAQEAJVCrj/9rQPDwJVCrj/9rQNDQJVCrj/+kALDAwCVQoECwsGVQq4//e0DAwGVQq4//hACg0NBlUKXRU7WRgrThD0KysrKysrKytd7U0QXV1x9isrKytN7QA/7T88MTABXSsAXQEzERQCBCMiJAI1ETMRFBYWMzI2EQRgwmT++9TO/vpwwketfda2Bbr8sd3+/KOOAQ3pA0/8sr+1YsIBFAAAAQAJAAAFRgW6AAoBPrECAkNUWEASBQEACAIBAgAICgAFCQgFAQIFL93NEN3NETMzAD8/PxESOTEwG0AkLwUBKgAoAyUKLwwwDGAMiQiJCZAMwAzwDAsgDFAMAgQCCwgCsQYCQ1RYtwkBDAsACAECAD8/ARESOTkbQCQKCQkgCAUUCAgFAAEBIAIFFAICBQkBAgXpIAoACAllCAFlAgi4/8BACyg5UAgBgAiQCAIIuAEBQA0CQCg5XwIBjwKfAgICuAEBQBEgBVAFAjAFYAWQBcAF8AUFBbgCiLMLYKgYKxkQ9F1x5F1xK+RdcSsYEO0Q7QA/PBoZ7Rg/PIcFLit9EMSHLhgrfRDEAUuwC1NLsBRRWliyAA8KuP/xsgkSAbj/8bIIFAK4/+44ODg4ODhZAUuwKFNLsDZRWli5AAD/wDhZWTEwAV1xXQBdWSEBMwEWFzY3ATMBAkH9yNIBfS4fIi0BjMb9wgW6+9eAcHh4BCn6RgAAAQAZAAAHdgW6ABgB20AmKQAmESkSJhg5ADYRORI2GEkARxFJEkcYWABXEVgSVxgQmAiYDwKxBgJDVFhAMxABGhkrFTQFNAxEBUQMSxVUBVQMWxVkBWQMaxV0BXQMexUPBRUMAwABEggACA8CCAIBAgA/Pz8/PxESFzldARESOTkbQB4DBAUFAgYHCAgFCgsMDAkNDg8PDBQTEhIVFhcYGBW4/zyzBQAYILj/PLMMEhEguP88QFoVCAkgAAUCAiABABQBAQAYBQgIHhUYFBUVGBIMCQkeFRIUFRUSEQwPDyAQERQQEBESCQwIGBUFDxEQDAACBRUMBQMYEA8PCQkICAICAQIYEhIREQAIGhcXGhBBCQFRACAADAFRABUBUQBAAAUBUbYgIAEBARkZuAGLsagYK04Q9F0aGU39Ghj9/RoZ/RhORWVE5gA/PBA8EDw/PBA8EDwQPBA8Ehc5ARI5ORESOTkREjk5ETk5h00uK4d9xIcuGCuHfcSHLhgrh33Ehy4YK4d9xCsrK4cOEMTEhw4QPMSHDhDExIcOEMTEhw4QxMSHDhDExAFLsA9TS7ARUVpYshIKGLj/9jg4WQFLsCVTS7AqUVpYuQAA/8A4WQBLsAtTS7AOUVpYswxABUA4OFlZMTABcl0hATMTFhc2NwEzExIXNjcTMwEjASYnBgcBAZ7+e8ffJBo4CgEX6tJPIxwt5sP+brv+yycHFxT+yQW6/D+XleskA979Gv7s84u0A676RgRdjCBlR/ujAAEACQAABUkFugATArVAKSYSARkBFgsCKRIpEzgBNwM4CDgJOA06DjUSNxMKEhMgEiE0EiASITQOuP/gsxIhNA24/+CzEiE0Cbj/4LMSITQIuP/gQGwSITQEIBIhNAMgEiE0dwF3CwImBCkHKAsqDiYSNgQ6CDoLOg41EkgIVARdCFwLWg5UEmcBZQRqCGsLaQ5lEnUEegh5C3oNdxJ3E4YEigeKCpUEuAi3EsYEyQjXBNgI2Q7WEucE6AjoDuYSLAa4/+pAEQwRAlUQFgwRAlULCAwRAlUBuP/4swwRAlWxBgJDVFhACwwAFRQQGAoRBlUGuP/oQA4KEQZVEAYAAg0ACAoCAgA/PD88ERI5OSsrARESOTkbQF0GBwgJCQEGBQQDAwsQEBMPDg0NARAQDRESExMLAQAJAg0LAwwTCgsBBhACEwkKExMgAAkUAAAJAwINDSAMAxQMDAMKCQkDAwICEw0NDAwACC8VARUXFxogDEAMAgy4AV+3IAqQCsAKAwq4Abi1XwKfAgICuAG4QAoGtEAQUBDPEAMQuAFfQAogABkUFcIhYKgYKytO9BoZTf1dGOUZ7V3tXf1dGE5FZUTmXQA/PBA8EDw/PBA8EDyHBU0uK4d9xIcuGCuHfcQAERI5OTk5Dw+HDhA8PAjEhw4QPDwIxIcOEDw8xIcOEMTExFkrKwArKzEwAV0AXQErKysrKysrK0NcWLkAC//eQAsZOQEiGTkOGBs5Erj/3rIbORO4/96yGzkEuP/oths5CCIbOQm4/8CyHDkNuP/AQB8cORNAHDkDQBw5DQ4WFzwTEhYXPQgJFhc8AwQWFz0LuP/eQC4SOQEiEjkLDB0hPQEAHSE8CwodIT0BAh0hPAsMExc9AQATFzwLChMXPQECExc8KysrKysrKysrKysrKysBKysrKysrKysrKytZAXEBXXEzAQEzARYXNjcBMwEBIwEmJwYHAQkCN/4M5wEKUyMxQwEn0/39Aivw/o8fITEV/pAC/AK+/oh1P1BXAYX9Tfz5AgstNVAe/gEAAAEABgAABUYFugAMAWq2CAk6AwQ7Cbj/57MSFzQIuP/nQA4SFzQEGRIXNAMZEhc0Cbj/2LMYITQIuP/YQDsYITQEKBghNBImBCkIKgovDgRoAWgGaAveBgQFBAMDBggHCQYGCQYDCQoMEAJVCSAKCxQKCgsGAwYJA7j/9kAWDBACVQMgAgEUAgIBBgwLBgEDAgABC7gCGUAJCgoJAwICAAgOuAIYQAkMCVJACoAKAgq4AbVADQsLDCAAA1JPAo8CAgK4AbVACQEBABQQEAJVALj/9kALDw8CVQAMDQ0CVQC4/+K0DAwCVQC4Ahi2DQ7CIWCoGCsr9isrKys8EPRd7RD9PBD0Xe0Q5gA/Pzw8PBD0PBESFzkBEjmHLisrCH0QxAWHLhgrKwh9EMSHDsTEhxAOxMRLsBdTS7AcUVpYtAgMCQwEuv/0AAP/9AE4ODg4WTEwAF0BXUNcWEAJCSIZOQgiGTkEuP/esRk5KysrWSsrKysrKysrKyERATMBFhc2NwEzARECO/3L7AEhUEVCXgEc4v23Am0DTf5GfHxzkAGv/LP9kwAAAQApAAAEsAW6AAwBDLESDrj/wEAPDRE0SAFHCEgJAwoICwkCsQYCQ1RYQA4MAA4NAQseDAgIBR4GAgA//Tw//cQBERI5ORtAK6sEAQMCAQEECQoECAoKJh0hNCgKAfkKAQogAQQUAQEECigLHDQBKAscNAi4/9izCxw0BLj/2EATCxw0AQoECAUeBwYCCwoeDAAICrsBtQABAAQBtUAbAAcwCEAIAghKDD8LAQsaDgEABQZRABkNtpkYK04Q9E30PBA8ThD2XTxN9HE8EOQQ/AA/PP08Pzz9PDwROQErKysrhwUuK11xK4d9xA4QxIcOEMTEAXJZMTABcV0rQ1xYQAkCIiE5ARghOQm4/961GTkCIhk5KysrK1kzNQE2NyE1IRUBByEVKQLvUEj8zgQa/MlZA6i0A6tkSq2t/AdnrQAB/+H+aQSK/usAAwAaQAwBPwACGgUAGQRDQRgrThDkEOYAL03tMTADNSEVHwSp/mmCggAAAgBK/+gEHAQ+ACgANwItQCwJDQkqGQ0aKikNKio5DTYVNxs6KkkqXQ1dKmoNaSpgMIoNhimaFpsaqQ0VKLj/6LQLCwZVJ7j/6EAZCwsGVaYZqii2GbsoxBnPKNIV3SgIRBYBHrj/9EARDAwGVRISDAwGVQUMDAwGVTW4/+BAVQwMBlUfFx8YKywqNDkEOSxJBEgsVghZK2YIaSt2DIcMyQz5DfkrETc0DgEEEC8kNBcyIRQYXylvKQIpHC8OPw6PDp8O/w4Fnw6vDu8OAw4MDw8CVQ64/+q0EBACVQ64//RAFRAQBlUODA0NBlUOBg8PBlUODhwDF7gCqrYYlRQcHAcAuP/0QBoMDAZVAEUnCjIcAwspYRBhAAYNDQJVACUhJLj/7LQQEAJVJLj/7EALDQ0CVSQEDAwCVSS4/+S0CwsCVSS4//S0CwsGVSS4/9xACxAQBlUkBg8PBlUkuP/8tAwMBlUkuAJbQA4nQAAmECYgJjAmryYFObj/wLQODgJVJrj/1rYODgJVJjE5uP/AQA0eIzQwOcA5AqA5ATkXuP/0QEEQEAZVFyUYIi8kvwbPBgIfBj8GAgYODw8CVQYMDQ0CVQYYDAwCVQYMCwsCVQYMCwsGVQYODQ0GVQYQDAwGVQYxOBD2KysrKysrK11x7fTtKxBdcSv2Kytd7fQrKysrKysrKzz9K+XlAD/tP+QrP+395BESOS8rKysrK11x7XEREjkREjk5ARESFzkxMABdKysrKwFxXSsrAHElBgYjIiY1NDY2NzY3Njc2NTQnJiMiBgcnPgIzMhYWFxYVFRQWFyMmAwYHDgIVFBYzMjY3NjUDPGS5aq+8R3NINWvaZwEzRYh/eR2wGG7QiYiqUBAJFyK8HBdixG9cMm1paKImHYNVRquFToFOFA4NGiQlCm4tPVlxGHGLS0BhSi548PuFPTgB3SgcEChNL0hgW089dwACAIb/6AQfBboAEAAdAYBAmwEFDA8kBTUFRQUFPx+wHwIfHyIcMxxCHHAfkB8GOhM8FjwaTBZMGl0IXQ1YD10WXhpqCGwNaA9uFm4awB/ZDNoX2hniE+wX7BnjHeAf/x8ZIAUvDy8UMAU/D0AFTA9QBWYF2h31BPoQDBAVDgQGAgAbHAYHAQoVHA4LGCTQCwEQC0ALYAuACwQfQA0NAlULDA8PAlULGA0NAlULuP/2tAwMAlULuP/wtAsLBlULuP/0tA8PBlULuP/gtAwMBlULuP/0QC8NDQZVC3QBETMABAwMAlUABA0NBlUAMwMlAgLAAQGQAaABsAHwAQQfAT8BTwEDAbj//rQQEAJVAbj//EAdDg4CVQEMDQ0CVQEQDAwCVQESCwsCVQEMCwsGVQG4//i0EBAGVQG4//xAFg8PBlUBGAwMBlUBFA0NBlUBGR5HNxgrThD0KysrKysrKysrK11xcjxNEP30KyvkEP0rKysrKysrK11x7QA/7T8/7T8RORESOTEwAF0BXXFyAHEhIxEzETYzMh4CFRAAIyInAxQXFjMyNjU0JiMiBgEtp7RysWKvcUD+8r28awI0VZF2rKV1dqwFuv31j0+PynP+7/7WnQGWv1WLzcvQxs0AAQBQ/+gD7QQ+ABoBWrECAkNUWEA0Dn8PAQ8LAUAAUABwAAMABBIcCwcYHAQLAQ4VBwgODgJVBwwNDQJVBwwMDAJVBxALCwJVBy8rKysrzdTGAD/tP+0QxF0yEMRdMjEwG0BHCQwBHxxDE0MXUxNTF2ATYBebApsDmg2kEKQaDAgNGQpqAmkDagV1DHANgA2mDLUJtgq1DAwWDIYM4wIDDiJfD28Pfw8DDwG4AqpAeTAAQABQAGAAcACQAKAA4ADwAAkADw8LAAAEEhwLBxgcBAscDwEPJA4IDQ0GVQ4iGwABACQLKx8BAQABAQFACwsGVQFAEBAGVQFIDAwGVQEaDQ0GVQFJHBUkzwcBHwc/BwIHDgsLBlUHChAQBlUHEgwMBlUHMRs0xBgrEPYrKytdce0Q9isrKytdcktTI0tRWli5AAH/wDhZ7XL0K+1yAD/tP+0SOS8ROS8QXeQQXeQxMABdcQFdcVkBFwYGIyIAETQSNjMyFhcHJiYjIgYVFBYzMjYDPLEd767a/vdy6Ymt3B+vGX9aiKqkhGqOAYUXt88BHQEKrAECga+hG2tsw9PWwoIAAAIARv/oA98FugARAB0BVUCkCgIEDSUNNA1EDQU1FDUcVwJUClIUUxxnAmQFZQljFGAcwB/UBdUT3RnlE+UU7xfrGeUd4B//HxYfHysaPBY8GksacB+QHwcuAiQNLhY6AjUNSwJFDUYUSRxXClYNZw3lBucW+gH0DhABFQMOCxAPABscCwcRAAoVHAMLGDMBACURDyUQENARARARQBFgEYARBB9ACwsCVR9ADQ0CVRESEBACVRG4//RAEQ8PAlURBg4OAlURGA0NAlURuP/yQAsLCwZVEQ4QEAZVEbj/7rQMDAZVEbj/+EBCDQ0GVRF0EiS/B88H3wf/BwQfBz8HTwcDBx4LCwJVBxgMDAJVBx4NDQJVBwwLCwZVBwwNDQZVBxoMDAZVBxkeNFAYK04Q9CsrKysrK11xTe39KysrKysrKysrK11xPBDtEP085AA/7T88P+0/PBE5ERI5MTAAXQFxXQBxITUGIyImJjU0EjYzMhYXETMRARQWMzI2NTQmIyIGAzhlxH/VdWrUg2CWL7P9IKx1dqWoe3ihhp6M+6OfAQOKUUECDvpGAhLMysHG2szEAAACAEv/6AQeBD4AFQAdAVNAFx8AHBUCVQNdBV0JVQtlA2sFbwllCwgVuP/ktA0NBlURuP/kQFINDQZVHRwNDQZVJxLZBfoU9hoEMRI6GTEcQRJNGkEcURJcGVIcYRJtGmEceAZ4FfYC9hgQABYBDw0XF1AWYBZwFgMWHA+QEKAQAhAQBBscCgcAugKqAAH/wLQQEAJVAbj/wEAQEBAGVRABAQGVExwECxdADbj/3LQNDQJVDbj/7rQNDQZVDbj/6rQMDAZVDbj/wEAJJyo0sA0BDRofuP/AsyUmNB+4/8BAQR4jNDAfAR8WMxAkB0AkKjQfBz8HTwcDByALCwJVBxgMDAJVBxwNDQJVBw4LCwZVBxwMDAZVBxYNDQZVBxkeNDcYK04Q9CsrKysrK10rTf3kThBxKyv2cSsrKytN7QA/7f1dKyvkP+0SOS9dPP1xPAEREjk5EjkxMAFdAF0rKysBcXIBFwYGIyIAERAAMzIAERQHIRYWMzI2ASEmJyYjIgYDXros7rnp/u8BFNzVAQ4B/OgKsoVjjP3aAlEMOFaJfKkBVhejtAEfAQMBDAEo/t7++RAgr7poAZWGQ2imAAEAEwAAAoAF0wAXAQ1AHhQJAQ8ZLxkwGUAZcBmbDJwNqQ0IGg0oDbAZwBkEGbj/wEAoGh80HQgNAwwPHAoBFQIrFBMEAwYACp8UART/E0AEFyUEAAMCkgEBALj/wLMxODQAuP/AQCscHzSQAAEZQA8PAlUZQA0OAlUAFBAQAlUAKA8PAlUAIg4OAlUALA0NAlUAuP/yQAsMDAJVABQLCwZVALj/6rQQEAZVALj/5rQPDwZVALj/+rcMDAZVAKMYGbwBugAhAPYBCgAYKyv2KysrKysrKysrKytdKys8EPQ8EDztEO3tXQA/Pzw8PP08P+05ETkxMEN5QBQQEQYJBwYIBgIGEAkSGwARBg8bASsBKyqBgQErcV0AcjMRIzUzNTQ3NjYzMhcHJiMiBhUVMxUjEbKfnxMag3ZMXBs4MlJEz88DmoxxazRGVxKdCkZgYoz8ZgACAEL+UQPqBD4AHgAqAW9AYAsLBRQsCyUUTAtFFAYJHRkdLAsmFCwjOQs2FEoLRhRWB1gLaAv6CvUVDi4jLCc+Iz4nTCeQLKAsBzYhNik/LEYLRiFFKVQhVClpB2MhYylgLIAs2ifoIe4j7ycRFxYGFbgCsbQoHBMHAbgCqkAQIAAwAGAAcACAAMAA0AAHALgCfUAyBRwcDwpFIhwMChYVMyUzCiUYGNAXARAXQBdgF4AXBCxACwwCVSxADQ0CVRcSEBACVRe4//RAEQ8PAlUXBg4OAlUXFg0NAlUXuP/qQAsLCwZVFxIQEAZVF7j/7rQMDAZVF7j//EBKDQ0GVRd0DwElACIfJL8Pzw/fD/8PBB8PPw9PDwMPIAsLAlUPGgwMAlUPIg0NAlUPHAsLBlUPDA0NBlUPGgwMBlUPGSssdCE0UBgrK070KysrKysrXXFN7fTtEP0rKysrKysrKysrXXE8EP3k9jwAP+3kP+39XeQ/7eQ/PDEwAV1xAF1xFxcWFxYzMjY3NicGIyICNTQSNjMyFzUzERQGBiMiJhMUFjMyNjU0JiMiBmavCzJDdH2IGA4BdrDb8G7Rjbx6pmXboL7qmaZ9fKitenioWBpRJTJkWjewiwE83ZgBAYyYgPxq+M94qwMq0cC/zMPGwwAAAQCHAAAD6AW6ABQBYbkAFv/AsxUXNAO4/+BADg0NBlUlBDUDRQO6DQQDuP/gQDoXGTQXCBEMERQDBQEADxwFBxQLCgwlCUAzNjT/CQHACQEWQAsLAlUWQBAQAlUJKBAQAlUJFA4OAlUJuP/sQBENDQJVCQQMDAJVCRoLCwJVCbj/9kALCwsGVQkUEBAGVQm4//hACw0NBlUJCg8PBlUJuP/2tgwMBlUJTha4/8BAFzQ2NLAW8BYCcBagFrAW/xYEFgIUJQEAuP/AQBAzNjTwAAEAACAA0ADgAAQAuP/6tBAQAlUAuP/6QBcODgJVAAQMDAJVAAgLCwJVAAQLCwZVALj/+kAWDw8GVQACDAwGVQACDQ0GVQBOFUdQGCsQ9isrKysrKysrXXErPP08EF1xK/QrKysrKysrKysrKytdcSvtAD88P+0/ETkROQESOTEwQ3lADgYOByUOBgwbAQ0IDxsBACsBKyuBACtdKwErMxEzETYzMhYWFREjETQmIyIGBhURh7R+wHauS7R1a1CNPAW6/fKSXaSc/V8CoYd7U459/bsAAgCIAAABPAW6AAMABwDNQF4JNgsLAlVPCZAJoAmwCcAJ3wnwCQcACR8JcAmACZ8JsAnACd8J4An/CQofCQEAAQcEAgMJBgN+AQAGBQYECgYHJQUABJ8EoASwBMAE4AQGwATwBAIABCAE0ATgBAQEuP/4tBAQAlUEuP/6QBcODgJVBAQMDAJVBAoLCwJVBBQLCwZVBLj/6rQQEAZVBLj//rQNDQZVBLj//EAKDAwGVQROCEdQGCsQ9isrKysrKysrXXFyPP08AD8/PD/tARESOTkREjk5MTABXXJxKxM1MxUDETMRiLS0tATrz8/7FQQm+9oAAAEAiAAAA/gFugALAmFAGwYMDQ0GVQcGVgZaCQMPDfMF9gYDCQwQEAJVBrj/9LQMDAJVCrj/9LQMDAJVCbj/9LQMDAJVA7j/6EAQDQ0GVVUDdwoCEgYgEyE0CLj/8LMSJzQJuP/wtBInNBIFuP/wsxIhNAm4//BAhBInNAYEBAUEBjcJRwQFJQYtClgKdwN1CtoD4wYHpgYBIwYmByUIOQY4CT8NTw1ZBFkGWAdZCX0EeQWZCcYG0gTWBuQG6Qf3BvkIFRIKCgUDAwQCBgYHCQkICgoFCQgIJQcGFAcHBgMEBCUFChQFBQoKCQYDBAgBAgAEBQYHCAgLCwAKBLgBD0AJBQQMDAZVBSIIuAEPQCEgBz8HAgcQDAwGVQcakA0BDQslAAIlAQGQAAE/AE8AAgC4//5AMQ4OAlUAEA0NAlUAEAwMAlUACgsLAlUAEgsLBlUAEgwMBlUACA0NBlUAGQwN4SFHZhgrK070KysrKysrK11xPE0Q7RDtThBx9itdTe30K+0APzwQPBA8Pzw/PBEXOYcFLisEfRDEhwUuGCsOfRDEBxAIPAg8AxAIPAg8sQYCQ1RYQA1LCQEfCYQDAgkYDRE0ACtdcVkxMAFDXFhACgksHTkJCB0dPAa4/96yHTkGuP/UsiA5Brj/1LEhOSsrKysrWV0AcV0BcQArK0NcWLkABv/AsiE5A7j/wLIWOQO4/96yEDkGuP/eshA5A7j/3rIMOQO4/96xCzkrKysrKytZASsrK0NcWEAS3QQBCBQWOQkIFBQ8CQgUFDwGuP/2shg5Brj/7LEbOSsrKysrAV1ZAF0rKysrKwFdcSszETMRATMBASMBBxGItAGq6f5qAb/e/qF/Bbr8vAGw/nb9ZAIfev5bAAABAIMAAAE3BboAAwDjtgU2CwsCVQW4/8CzNzg0Bbj/wLM0NTQFuP/AszAxNAW4/8CzIiU0Bbj/wEAlFRc0DwUfBZ8F3wUETwXfBfAFAx8FcAWABf8FBAEAAAoCAyUBALj/wLM3ODQAuP/AQBUzNTSfAAHAAPAAAgAAIADQAOAABAC4//i0EBACVQC4//pAHQ4OAlUABAwMAlUACgsLAlUAFAsLBlUACBAQBlUAuP/+tA0NBlUAuP//tAwMBlUAuP/8QAoMDAZVAE4ER1AYKxD2KysrKysrKysrXXFyKys8/TwAPz8xMAFdcXIrKysrKyszETMRg7QFuvpGAAABAIcAAAYmBD4AIwHHuQAN//S0DQ0GVQi4//S0DQ0GVQm4/9hATQsNNCUE5ATkCeEX5SAF1QX2IAIXCCAjCRgbIAkDAyMeHAYVHAsLBgcBBiMaGRAK0CUBkCWgJQIlFxcaDiWQEQERBBAQAlURGA8PAlURuP/sQAsODgJVERQMDAJVEbj/6EAXCwsCVRECCwsGVREMEBAGVREGDw8GVRG4//q0DAwGVRG4//i0DQ0GVRG4AV1ADBglkBsBGxgPDwJVG7j/7EALDg4CVRsUDAwCVRu4/+5AEQsLAlUbBAsLBlUbChAQBlUbuP/+QAsNDQZVGwwPDwZVG7j//LQMDAZVG7gBXUAWAAIzIyUB0AABkACgAAIfAD8ATwADALj//kAdDg4CVQAQDQ0CVQAQDAwCVQAMCwsCVQAWCwsGVQC4//y0EBAGVQC4//RAFA8PBlUACgwMBlUADg0NBlUAGSQluAF4syFHUBgrK070KysrKysrKysrXXFyPE395BD0KysrKysrKysrXe30KysrKysrKysrK139TkVlROZxcgA/PDw8Pz88TRDtEO0RFzkBERI5EjkxMEN5QA4MFBMmFAwRGwESDRUbAQArASsrgQFdAF0rKyszETMVNjYzMhYXNjMyFhURIxE0JiYjIgYVESMRNCYjIgYGFRGHoTKmanaXH37KnqqzI1w+cJS0WGRMgToEJpVOX2JYuq+2/ScCnWxfOpWk/ZcCsnh4UJqR/dkAAAEAhwAAA+YEPgAWAX1AEwUDBhMCqBC4EOMD5xPwA/YTBgS4//BAPAsNNHkQAZgQ0BjgGP8YBCAIFA4UFhIcBQcBBhYNCg0ODA4kGEAQEAJVGEALCwJVCygQEAJVCxQODgJVC7j/7EARDQ0CVQsEDAwCVQsiCwsCVQu4//RACwsLBlULFBAQBlULuP/5QAsNDQZVCwoPDwZVC7j/9kASDAwGVQtAMzY0/wsB/wsBC04YuP/AQBo0NjSwGPAYAnAYoBiwGMAYBBgDAjMVFiUBALj/9rQREQJVALj/+rQQEAJVALj/+kAXDg4CVQAEDAwCVQAKCwsCVQAECwsGVQC4//pAEQ8PBlUAAgwMBlUABA0NBlUAuP/AQBIzNjTwAAEAACAA0ADgAAQAThcQ9l1xKysrKysrKysrKzz9PPQ8EF1xK/ZdcSsrKysrKysrKysrKyvtPBA8AD88Pz/tETkBEjkxMEN5QBYGEQkKCAoHCgMGECYRBg4bAQ8KEhsBACsBKysqgQFdcQArXXEzETMVNjMyFhYXFhURIxE0JiYjIgYVEYeidd1goVAQCrQqa0hzpwQml69FcE0yff1zAoZubUGSzP28AAACAET/6AQnBD4ADQAZAWu2FRgNDQZVE7j/6LQNDQZVD7j/6EBzDQ0GVRkYDQ0GVRIHChkMRwZICFYGWQhnBmkICDQQOhI6FjUYRRBLEksWRRhcBVwJUhBdEl0WUhhtBW0JZBBtEm0WZBh3ARUJBgUNWwNUBVQKWwxsA2UFZQpsDAoXHAQHERwLCxQkG0ANDQJVG0ALCwJVB7j/6kARDw8CVQcYDQ0CVQcQCwsCVQe4//C0CwsGVQe4//C0DQ0GVQe4//C0Dw8GVQe4//C0DAwGVQe4/8BAEyQlNDAHAQAHEAcgBwMHMd8bARu4/8BASR4jNDAbARsOJAAMDg8CVQASDQ0CVQAMDAwCVQAcCwsCVQAOCwsGVQAODQ0GVQAMEBAGVQAWDAwGVQBAJCU0HwA/AAIAMRo0NxgrEPZdKysrKysrKysr7RBxK132XV0rKysrKysrKysr7QA/7T/tMTABcV0AcUNcWEAJUwVTCWIFYgkEAV1ZACsrKysTEDc2MzIAFRQGBiMiABMUFjMyNjU0JiMiBkSkicXbARZ764vf/u25soeGsrOFh7ICEwEnjnb+4f3N64IBHgENzMvM0cXLygACAIf+aQQhBD4AEgAeAWJAjgwQLRA9EEsQBD8gsCACHyApDCMdMhUyHUIdcCCQIAg6FzobShdKG1kIWwxcF1wbaghrDGkQbRdrG8Ag0xTdGN0a0x7kFOQe4CD/IBYjBCsQKxU1BDoQRgRKEFoQ5QvrHf4QCxEOAxYcHAYHAQYWHA4LAA4ZJNAKARAKQApgCoAKBCBACwsCVSBADQ0CVQq4/+ZACw8PAlUKGA0NAlUKuP/6tAwMAlUKuP/utAsLBlUKuP/0tA8PBlUKuP/oQCMMDAZVCnQBEzMCMxIlAADAAQGQAaABsAHwAQQfAT8BTwEDAbj//EAdDg4CVQEQDQ0CVQEQDAwCVQEQCwsCVQEMCwsGVQG4//a0EBAGVQG4//xAFg8PBlUBDAwMBlUBEg0NBlUBGR9HNxgBK04Q9CsrKysrKysrK11xcjxNEP305BD9KysrKysrKytdce0APz/tPz/tETkSOTEwAF0BXXFyAHETETMVNjYzMhYWFRQCBiMiJicRAxQWMzI2NTQmIyIGh6Q6kmiI0Gp133tajy4RpnZ4q6d0c7H+aQW9ilFRjP+Yo/77i0w6/fsDpM3Ey9XLytcAAAIASP5pA+AEPgAQABwBNkCOCwIrAioYOwJLAnkMBj8VPxlLGZAeoB4FNBM0Gz8eRBNEG1MTUxtjE2MbYB6AHtQG1RLmBukM6hgQKQIiDCsVOQI1DEkCRgxaAmkC2QzbGOMW6RnmG/wCDwEEDRQaHAsHDgYUHAQLAA4XDjMAJRAQ0A8BEA9AD2APgA8EHkALDAJVHkANDQJVDxIQEAJVD7j/9EARDw8CVQ8GDg4CVQ8WDQ0CVQ+4//5ACwwMAlUPFhAQBlUPuP/otAwMBlUPuP/0QD8NDQZVD3QRJL8HzwffB/8HBB8HPwdPBwMHJAsLAlUHGgwMAlUHIg0NAlUHFgwMBlUHGg0NBlUHGR0edCE0UBgrK070KysrKytdcU3t/SsrKysrKysrKytdcTwQ/fQ8AD8/7T8/7RE5EjkxMABdAV1xAHEBEQYGIyIAETQ2NjMyFzUzEQEUFjMyNjU0JiMiBgMsKpdVvf7vb9N+xXGi/SGseHOmr3Z1o/5pAgg7TgEuAQeg/oOmjvpDA63NzcPH1NbHAAABAIUAAALGBD4AEQDJQDsvEwEQBAEjBDQEQwRTBGYEdAQGCREICQgJDRMRCQ0AAwgBCxwGBwEGAAoJKJAIAQgiIBMBEwIiESUBALj/wEAQMzY08AABAAAgANAA4AAEALj/+LQQEAJVALj/+EARDg4CVQAEDAwCVQAGCwsCVQC4//y0EBAGVQC4//RAFg8PBlUABgwMBlUACA0NBlUAThJHxBgrEPYrKysrKysrK11xKzz95BBd9HLkAD8/P+0ROTkROTkBERI5OQAQyYcOfcQxMABdcgFdMxEzFTY2MzIXByYjIgYHBhURhaI+aT9bXj5CQjteFB4EJqFxSDqnJ0c/YHL91AAAAQA//+gDsQQ+ADADF0B7BCIUIjoJSglEJFYiZSJ8CY4JhCSmE6sswgMNCRcaGBcwSyzWFwUbAlUCAhAyAQoYXAhcCVwKXAtcDFwNaghqCWoKagtqDGoNtCa0Jw8nJiQnJCk2JFoKWQtkJmQodCN0JIAkkwqcDJIolyyVMKQKqQyjJ6QosybFJhYouP/0tA0NBlUiuP/0tA0NBlUjuP/0tA0NBlUkuP/0tA0NBlUouP/0tAwMBlUiuP/0tAwMBlUjuP/0tAwMBlUkuP/0tAwMBlUduP/eQBIeOVoIJyUMCgQaICYVBAsuHRq4AqpAIhksCwsCVR8ZPxlPGV8ZrxnPGQYPGR8ZbxnfGQQfGY8ZAhm9AlUAFQAAAqoAAf/AQBQLCwJVEAFAAQIQAdABAgABEAECAbj/wLMUFjQBuP/AQBAOETQBAS5cHWwdAh0cFQcEuP/0tAsLAlUEuP/mtBAQBlUEuP/mQBMPDwZVBBwuCx8aARokGUATGDQyuP/AQC8PDwJVGRgPDwJVGRgNDQJVGRYMDAJVGSAQEAZVGSAPDwZVGRAMDAZVGRYNDQZVGbgCW7IHJCq4/8C1HDnQKgEquP/mtAwMAlUquP/otA8PAlUquP/otAwMBlUquP/qtg0NBlUqGjK4/8BAIScqNGAywDICPzKAMgIyEAEBASQAGA0NAlUAEA0NBlUAILj/9LQNDQJVILj/9LQQEAZVILj/9EAZDw8GVSAkDxALCwJVDxYMDAJVDyANDQJVD7j/+kAgDw8CVQ8ODAwGVQ8MDQ0GVQ8i3wABPwBPAAIAGTE0NxgrThD0XXFN9CsrKysrK+0rKysQKyvtck4QXXEr9isrKytxK03t9CsrKysrKysrK+1yAD/tKysrP+1xEjkvKytdcXIr5BD9XXFyK+QREjkREjkBERIXOTEwQ3lAQCctHiMFFCwmERASEBMQAwYiDSAbAAkoBxsBBS0HGwEeFCAbACEOIxsAIiMNDAgpChsBKCcJCgYrBBsAHxAdGwEAKysQPBA8KxA8EDwrASsrKysqK4GBgQArKysrKysrKytdcQFdcnFdEzcWFjMyNjU0JyYnLgI1NDY3NjYzMhYWFwcmJiMiBhUUFxYXFhceAhUUBgYjIiY/sg+Je3x4NSWTxplPQTgqkVN9vVoRsAxzaXxqFhYvG4S/l1Zpxn3P2QE9HGtyZUQ9IxglMkmBTkd5KB8rSHtnGFJcUjcjHB0TCiQzQXxcWp9XrAAAAQAk//ICKgWZABcA2LkACv/AsyMmNAm4/8BAQSMmNIAZAQABDA0KAQMAFhAJKw8KBhYcAwsPECIAIgENEiUMAf8HCEUJRWAHcAeAB5AHBAAHIAegB7AHwAfQBwYHuP/utBAQAlUHuP/0tA8PAlUHuP/ytA4OAlUHuP/4tA0NAlUHuP/4tAwMAlUHuP/6tBAQBlUHuP/wQAsPDwZVBwYMDAZVB7j/6LQNDQZVB7oCagAYATaxZhgrEPYrKysrKysrKytdcfTkEO08/TwQ5PQ8AD/tPzz9PBE5EjkRMzMQyTEwAV0rKyUXBiMiJiY1ESM1MxE3ETMVIxEUFhYzMgIQGkw8YmwshISztbUTKygeoZ8QPmWiAmOMAQds/o2M/ZNNLBoAAAEAg//oA+AEJgAYAU+5ABr/wEAJFRc0AiATFjQPuP/wQDMSFDQrEwEkCBMWDAETFgsGAAoRHAMLADMWJRgXQDM2NBpAEBACVRcoEBACVRcSDg4CVRe4/+xACw0NAlUXBAwMAlUXuP/0QAsLCwZVFxQQEAZVF7j/+EALDQ0GVRcMDw8GVRe4//ZADQwMBlX/FwHAFwEXThq4/8BAFTQ2NLAa8BoCcBqgGrAa/xoEGgwlCbj/wEAQMzY08AkBAAkgCdAJ4AkECbj/+LQQEAJVCbj/+EARDg4CVQkEDAwCVQkKCwsGVQm4//ZAFg8PBlUJAgwMBlUJAg0NBlUJThlHUBgrEPYrKysrKysrXXEr7RBdcSv2XXErKysrKysrKysrKzz95AA/7T8/PDk5ARESOTEwQ3lAGgQQDg0PDQIGBwgGCAUIAwYQBAwbAA0IERsAACsBKyoqgQBdASsrKyE1BiMiJiYnJjURMxEUFxYWMzI2NjURMxEDP3zVXqNPEAu0CxFuUVGOO7SctEhtTzVzApL9s40xR1FTj4gCOfvaAAEAGgAAA+gEJgAKAeqxAgJDVFhAFwUIAAoIBgEGCgAFCQgFAQIFJA8PAlUFLyvdzRDdzREzMwA/Pz8SOTEwG7c1BQEAIhE5Crj/3kANETkJFhIcNAgWEhw0Arj/6rMSHDQBuP/qsxIcNAq4/9hACR4hNAAoHiE0Crj/6EAJIiU0ABYiJTQKuP/aQH4oLjQAICguNA8MKQAoCSYKOQA1CkgARwpWAVYCWQhYCWYBZgJpCGkJeAB3AXcCeQh4CXcKhwGHAoYDiQeICIoJnQCYCZEKrACiCr0AtwexCskAxQraANUK7ADjCvsA9AosCgAFChgAFgooACYKNwpPAEAKCQVAEhY0BUALDTSxBgJDVFhACQUBAAgGAQYACrj/9EAPDQ0GVQoADA0NBlUABQkIuP/0QBINDQZVCAUBAgwNDQZVAgUFDAsREjkv3SvNEN0rzRDNK80rAC8/PxESOTEwG0A3CgcICCUJChQJCQoAAwICJQEAFAEBAAUKCgAKCQgIAgIBBgcKCQMAAQUvDAEMIghAQEAJgAkCCbgBG7VABYAFAgW4ARtACSACQAEiC+rSGCsQ9u0aGf1d/V0aGO3kXRESOTkSOTkAPzwQPBA8PzwROYcFLiuHfcSHLhgrh33EWTEwACsrAXFdKysrKysrKysrKysrAF1ZIQEzExYXNjcTMwEBrv5svuQlHxgr7Ln+bgQm/YRnb1R2Aoj72gAAAQAGAAAFtwQmABIEHbECAkNUWLkAEv/0QBENDQJVBwYNDQJVAAYNDQJVCrj/1LQMDQJVBLj/6EALDA0CVREgDA0CVQq4/8C0DhACVQS4/8BALw4QAlURQA4QAlUEChEDAQAMBgcGAQYPCgAKDQwGDAwCVQwRAQIECgQRCgwMAlURuP/4tA0NAlURLysrzc0Q1s0Q1CvNAD8/Pz8/ERIXOTEwACsrKysrKwErKysbQBYPFAEqBCkKAkoRWxGOEQMRIA0NBlUKuP/gtA0NBlUEuP/gtA0NBlURuP/wQAkfITQQHB0nNAm4//BAtx8kNAQGDAkTBhsJGRIFBAAEBgsJCw4IEhAAEwMUBxwIGwsdDiQAJQcqCCsONAA1BzoIOw5EA0cGQAdNCEsLQw9HEUoSWw9SEmsHZAhnEnkGegd0CLkGug+2EvUG+wkoCxEoACgNJw4oDycSLxQ4ADcSdwiGCJgDlwynAagCqAumDLUAtga6DsgE1gbZCegE6A/nEvQG+gkcCwYNDQZVDAYNDQZVEAYNDQZVDgYNDQZVDwYNDQZVErEGAkNUWEAbCg4PBBIAEQgHCCUHDyUOEiUAAA4HAw0BDCUNuP/WQDcLCwZVDQIlASoLCwZVAQ0BFBMGCgsRJgorEVQEUgpcEWwRfBGKEQoRCgQDAAEPCgAKDAYHBgEGAD8/Pz8/ERIXOV0BERI5OS8r9C8r9BESFzkQ5BDkEOQREjkREjkREjkbQBQDBQUCBgcHBQkKCggLDAwKEBERD7j/S7MFABIguP9JQGYKDw4gwxEHCCAHERISKwUHFAUFBw4KDAwlDQ4UDQ0OCBEPDysKCBQKCggABQICJQEAFAEBAAACAQcSBAgPEQwODQoRCgQDEg0MDAgIBwcCAgEGEg8PDg4AChT2EA0BYA1wDYANAw24AadACiBPCgFvCn8KAgq4AlVACU8RAW8RfxECEbgCVUALEAUBYAVwBYAFAwW4Aae1AfYT9mYYK04Q9BlN9F1dGP1dcf1dcRoZ/V1dGOYAPzwQPBA8PzwQPBA8EDwQPBIXOQEREjk5Ejk5ETk5Ejk5h00uK4d9xIcuGCuHfcSHLhgrh33Ehy4YK4d9xCsrK4cOEMQHDhA8Bw4QPIcOEMSHDhDES7AfU1i0DSAMIAK8/+AAAf/gAA7/0LQAMA8gErj/4AE4ODg4ODg4OFlLsDRTWLkACP/QsQcwATg4WUuwIVNLsDNRWli5AAj/4LEHIAE4OFlLsBJTS7AeUVpYuQAO/9C2DyANIAwgCLj/0LIHMBK4/+CyADgCuv/gAAH/4AE4ODg4ODg4ODg4WUuwElNLsBdRWli5ABH/4LMKIAQgADg4OFlZMTABQ1xYuQAO/9S2EjkALBI5ALj/1LETOSsrK1krKysrK11xcisrKwArKytxXQFdWSEBMxMXNjcTMxMXNxMzASMDJwMBS/67uqk/BDOpuZ81Pbav/rS7qSnXBCb9m+QRygJu/ZjLzQJm+9oCfLX8zwABAA8AAAPxBCYAEAHcsQICQ1RYQBUPAQsGBAIJBgIGDQoACg8YDw8CVQ8vKwA/Pz8/ERc5MTAbtw8SAQ8iGTkGuP/eQFAZOVoPlgSWCJkOmg/ABcAGwAfLDwkPQBY5GgMTCRUNGhA1AToLgQGOCwgvElcEWQdZC1gOlwGYCpgLtwK4DMgLyg7MENoD1QnRDdsQ5QoSErEGAkNUWEALDAASEQ8YDRAGVQa4/+hADg0QBlUPBgACDQAKCgIGAD88PzwREjk5KysBERI5ORtAZgYGAwcICQkBBgYJBQQDAwsPDxAODQ0BDw8NEAsBAAkCDQsDDBAKBg8CDwoQxgDGCQIQJQAJFAAACQMCDcYNAQ0lDAMUDAwDCgkJAwMCBhANDQwMAApPEgESSQ1+DCIKD2EGCX5ACrgBG7dABlAGgAYDBrgCQ0AOIAN+AiJPAAEASRF8xBgrEPZd9O0aGf1d/RoY7RDlEPTt5l0APzwQPBA8PzwQPBA8hwUuK12HfcSHLhgrXX0QxAAREjk5Dw+HCMSHDhDECMSHDhDExAjEBw4QPDwIPFkxMAFDXFi0DhgdOQu4/95ACx05DCIXOQMiFzkLuP/esiE5ELj/wEAKFTkBIiE5CUAcOSsrKysrKysrWV1xACtdKysBXVkzAQEzFxYXNjc3MwEBIwMnAQ8BhP6Z4aMuHCwls9f+kQGL3do6/ukCKAH++UcwQjP7/gz9zgFKWf5dAAEAIf5RA+4EJgAaAfexAgJDVFhAHQoUDwMLAxwZDxIGCwYTQBIPIAtADCAPGA8PAlUPGS8rGt0aGM0aGRDdGhjNAD8/P+0SFzkxMBuzDxwBD7j/3kBtHDkoFFYPrwoDQA1ADwIPICgwNBAgKDA0BwwJEhYNGBInCycMJw02DDYNNQ6ZEQsoEigTSBZZElkTWRVpEmkTaRV5BnYNeRF6FHoVhQ2KEYwSjBOJFJgKqAu8ELsRuhTqCucU9Q39EPkU/xweErEGAkNUWEAWEwscGwQPRA+EDwMPGQsDHBkPEgYLBgA/Pz/tERI5XQEREjk5G0A3Dw8MEBESEgoAAxkUExMlEgoUEhIKDwwPEQwlCwoUCwsKExISDAwLBgMcGQ8AHBAcAi8cvxwCHLgCP7UPE0ASQBS4AlRACz8SQBICXxK/EgISuAFCtg8BIgBFGwq4AlRAEg8gC0BAIAwwDE8MA1AM/wwCDLgBQrMvDwEPuAI/tBsgfGYYKxoZEP1x9F1xGhjtGhkQ7RgQ9OQZEORdce0aGBDtGRDkXXEAGD/tPzwQPBA8hwUuKwh9EMSHBS4YKw59EMQAERI5hw4QPDwIxEuwDlNLsBhRWli7AAz/6AAL/+gBODhZWTEwAUNcWLkAFP/etjc5CiI3OQ64/+i1FTkRIhU5KysrK1ldcSsrAHFdKwFdWRMnFjMyNjc2NzY3ATMTFhc2NxMzAQYHBgYjIn8UOyw8SBcRJgUL/m3C3SsiHyvjtP5sQSQwfFY0/mepECgkG2sPHQQo/Zl1gXx2Amv7yK9CWVMAAAEAKAAAA9QEJgAOAa9ADRK4AskIAhIBMhIXNAi4/85ACRIXNAE+HiE0CLj/wkBKHiE0KQIoCS8QOQE5CkkBRgJGCEkJTxBcAVQCVAhaCVAQbAFjAmMIagl7AXQIewmLAYUIiQn5AfQCGxkIJgEpCCsJOQilCNcBBxC4/8C3EBU0AiwSOQm4/9RAIxI5AQI6CQoCCAoKJQECFAEBAgENDggGAmEFKwcGBgphDQANuP/0QAkLCwZVDSsOCgK4AQ+0CAgHBQa7AlsAAAAH//RAFgsLBlUHIg2gDgEADkAOYA6ADvAOBQ64//RAJAsLBlUOdAAKfgEBrwABTwBvAP8AAwAYCwsGVQAZDxB0IXzEGCsrTvQrXXE8TRDtEP0rXXE85CsQ9DwQPBD9AD/tKzwQ5T88/eURORESOYcFLiuHfcQQDsQrMTABKysrcV0AKysrK0NcWLUpASYIAgG4/85ACRIXNAgyEhc0Abj/wrceITQIPh4hNAArKysrAXFZAV1DXFi5AAj/3rIPOQm4/96yDzkJuP/otxs5CQgWGz0JuP/wshc5Cbj/+EAKFjkCFBY5AhoWOSsrKysrKysrWTM1AQYjITUhFQEHNjMhFSgCpHNY/k8DZP3Bb3lqAeuSAwgGknf9XnsJmwAAAwAD/+4F6AXTAA8AHwA6ATNAIJQSlBabGpsepgOoC6gNuTDUEtQW2xrbHtUz1jYOcAgguAKrsyGHJC+4AquzMC4BLrsCYAArADgCYkAQTyQBDyRvJH8k7yQEJJQIMrgCYkALACuPK/8rAyuUABi4AmKyCAsQuAJisgADL7gCYrIu0yC4AmKzIYgENb0CYgAnAmQADAAcAmKzBBo8FLgCYrUMGTuzehgrThD0Te1OEPZN7RD07RD07fTtAD/tP+0Q9F3tEPRdce0Q/V3kEP3kMTBDeUBUMzclKgEfKSYSJQ4mAiUeJhYmCiUGJholMyo1HwA3JTUfABEPFCEAHwEcIQEXCRQhABkHHCEBNCgyHwE2JjgfABMNECEBHQMQIQEVCxghABsFGCEAKysrKysrASsrKysrKysrKysrKysrK4GBgQFdATIEEhUUAgQjIiQCNTQSJBciBAIVFBIEMzIkEjU0AiQTFwYGIyImNTQ2NjMyFhcHJiYjIgYVFBYzMjYC9r4BasrH/pnExP6ZyMsBar6f/tOqpwEso6MBLKap/tJUex7Di7DcZLl3hbAgdx51T3OVjXBaiAXTw/6VxcP+mMfHAWjDxQFrw32j/tGko/7Vp6cBK6OkAS+j/RAkfZXkyoTDY39tHUpPpJmZnWgAAAH//AHKBG8CWwADAB5ADwE1AAIaBSAAAQAZBLN6GCtOEORdEOYAL03tMTADNSEVBARzAcqRkQAAAQAAAAU4UgAAAABfDzz1CDsIAAAAAACi4ycqAAAAANKUfxr6r/1nEAAIDAAAAAkAAQABAAAAAAABAAAHPv5OAEMQAPqv+noQAAABAAAAAAAAAAAAAAAAAAANXQYAAQAAAAAAAjkAAAI5AAACOQCwAtcAXgRzABUEcwBJBx0AdwVWAFgBhwBaAqoAfAKqAHwDHQBABKwAcgI5AKoCqgBBAjkAugI5AAAEcwBVBHMA3wRzADwEcwBWBHMAGgRzAFUEcwBNBHMAYQRzAFMEcwBVAjkAuQI5AKoErABwBKwAcgSsAHAEcwBaCB8AbwVW//0FVgCWBccAZgXHAJ4FVgCiBOMAqAY5AG0FxwCkAjkAvwQAADcFVgCWBHMAlgaqAJgFxwCcBjkAYwVWAJ4GOQBYBccAoQVWAFwE4wAwBccAoQVWAAkHjQAZBVYACQVWAAYE4wApAjkAiwI5AAACOQAnA8EANgRz/+ECqgBZBHMASgRzAIYEAABQBHMARgRzAEsCOQATBHMAQgRzAIcBxwCIAcf/ogQAAIgBxwCDBqoAhwRzAIcEcwBEBHMAhwRzAEgCqgCFBAAAPwI5ACQEcwCDBAAAGgXHAAYEAAAPBAAAIQQAACgCrAA5AhQAvAKsAC8ErABXBVb//QVW//0FxwBoBVYAogXHAJwGOQBjBccAoQRzAEoEcwBKBHMASgRzAEoEcwBKBHMASgQAAFAEcwBLBHMASwRzAEsEcwBLAjkAvQI5ACMCOf/lAjkACQRzAIcEcwBEBHMARARzAEQEcwBEBHMARARzAIMEcwCDBHMAgwRzAIMEcwBJAzMAgARzAGsEcwAbBHMAUQLNAG0ETAABBOMAmQXlAAMF5QADCAAA4QKqAN4CqgA9BGQATggAAAEGOQBTBbQAmgRkAE4EZABNBGQATQRz//0EnACgA/QAOAW0AHoGlgChBGQAAAIxAAAC9gAvAuwALQYlAH8HHQBEBOMAgQTjAJ4CqgDoBKwAcgRkAFQEcwAuBGQAMwTlABoEcwCGBHMAjAgAAO8FVv/9BVb//QY5AGMIAACBB40AUgRz//wIAAAAAqoAUwKqAEcBxwCAAccAbARkAE4D9AAvBAAAIQVWAAYBVv45BHP/5AKqAFwCqgBcBAAAFwQAABcEcwBJAjkAuQHHAGwCqgBHCAAAJQVW//0FVgCiBVb//QVWAKIFVgCiAjkAjQI5/+ACOQAEAjkAFQY5AGMGOQBjBjkAYwXHAKEFxwChBccAoQI5AMYCqgAZAqoABgKqAB0CqgAuAqoA5QKqAKICqgBrAqoAOgKqAEsCqgAoBHMAAAHHAAMFVgBcBAAAPwTjACkEAAAoAhQAvAXH//0EcwBJBVYABgQAACEFVgCeBHMAhwSsAHIErAChAqoAawKqABkCqgAhBqwAawasAGsGrAAhBHMAAAY5AG0EcwBCAjkAsQVWAFwEAAA/BccAZgQAAFAFxwBmBAAAUARzAEYEa//hAqoA7gVW//0EcwBKBVb//QRzAEoFxwCeBOsARwXH//0FVgCiBHMASwVWAKIEcwBLBHMAlgHHAEIEcwCWAlUAiARzAJoCrACDBccAnARzAIcFxwCcBHMAhwY5AGMEcwBEBccAoQKqAIUFxwChAqoAPAVWAFwEAAA/BOMAMAI5ACQE4wAwAwAAIwXHAKEEcwCDBccAoQRzAIME4wApBAAAKATjACkEAAAoBGgApAY5AGAGYgBVBKAASAR0AEgDkQBiBPAARAMpAC4FMABIBGv/4QQAALAC6wBSCMAAMwgAAE8EAACZCAAATwQAAJkIAABPBAAAmAQAAJgH1QFqBcAAngSrAHIE1QCdBKwAcQTVAiIE1QEFBav/6QUAAckFqwJ+Bav/6QWrAn4Fq//pBasCfgWr/+kFq//pBav/6QWr/+kFq//pBasBwAWrAn4FqwHABasBwAWr/+kFq//pBav/6QWrAn4FqwHABasBwAWr/+kFq//pBav/6QWrAn4FqwHABasBwAWr/+kFq//pBav/6QWr/+kFq//pBav/6QWr/+kFq//pBav/6QWr/+kFq//pBav/6QWr/+kFq//pBav/6QWr/+kFqwLWBasAZgWr/+oF1f//BNUAkggAAAAH6wEwB+sBIAfrATAH6wEgBNUAsgTVAIAE1QAqCCsBmAhrAbgHVQAQBgAA9AYAAG8EQAA6BUAANwTAAD8EFQBABAAAJQYAAFUF4QC/A40AiQTV/9kBgACAAtUAhgcVAGEClgAPBNUAkgLWAIMC1gCDBNUAsgLWAHAFVv/9BHMASgXHAGYEAABQBccAZgQAAFAFVgCiBHMASwVWAKIEcwBLBVYAogRzAEsGOQBtBHMAQgY5AG0EcwBCBjkAbQRzAEIFxwCkBHMAhwXHAB8EcwAGAjn/zgI5/84COf/kAjn/5AI5//YCOf/1AjkASwHHABkEAAA3Acf/ogVWAJYEAACIBAAAhgRzAJYBx//6BccAnARzAIcFyQClBHMAiwY5AGMEcwBEBjkAYwRzAEQFxwChAqoAawVWAFwEAAA/BOMAMAI5AAwFxwChBHMAgwXHAKEEcwCDBccAoQRzAIMFxwChBHMAgweNABkFxwAGBVYABgQAACEBxwCJBVb//QRzAEoIAAABBx0ARAY5AFME4wCBAjkAuQeNABkFxwAGB40AGQXHAAYHjQAZBccABgVWAAYEAAAhAccAigKq/+EEcwAbBM0AWgasAGsGrAAiBqwAIgasAEoCqgDiAqoAawKqAN4Cqv/qBVf//wZG/6cGtP+oAxL/qAYy/6cG2P+nBgX/pwHH/3gFVv/9BVYAlgVY//4FVgCiBOMAKQXHAKQCOQC/BVYAlgVYAAsGqgCYBccAnAUzAG0GOQBjBccApAVWAJ4E8gCUBOMAMAVWAAYFVgAJBq8AfwX7AGECOQAEBVYABgSgAEgDkQBiBHMAiwHHAGsEYACIBJoAjAQAABkDhwBIBHMAiwRzAFwBxwCJBAAAhgQAABgEnACgBAAAGgOVAFwEcwBEBI0AgwPbAFYEYACIBDMAEQW0AHoGPwBXAcf/yQRgAIgEcwBIBGAAiAY/AFcFVwCiBusAMgRVAKEFwABkBVYAXAI5AL8COQAEBAAANwh1AA0IFQCkBtUAMQSpAKEFFQAKBcAAoAVW//0FQACnBVYAlgRVAKEFawAABVYAogdjAAcE1QBOBcAAoQXAAKEEqQChBUAAEgaqAJgFxwCkBjkAYwXAAKAFVgCeBccAZgTjADAFFQAKBhUAUgVWAAkF6wCfBVUAVwdVAKEHgAChBlUAAAcVAKgFQAClBcAAVQgVAKQFxwAaBHMASgSVAFsEQACIAusAiASrAAAEcwBLBVr/+wOrADIEeACHBHgAhwOAAIYEqwAYBYAAjARrAIgEcwBEBFUAiARzAIcEAABQA6oAJgQAACEGlQBLBAAADwSVAIoEKwBFBmsAjQaVAI0FAAAoBcAAiwQrAIQEFQAwBgAAiQRVAB8EcwBLBHMAAALrAIkEFQBLBAAAPwHHAIgCOQAJAcf/ogdAABMGgACDBHMAAAOAAIYEAAAhBGsAiAPpAKEDSgCICAAAQQiVAKAFhQAtAAABAQAAAB4AAAAxAAAAMQAAAQEAAAB+AAAAfgAAAIwAAACMAAABAQAAABAAAAEBAAABIQMQAH0AAACMAjMA0gAAAwsAAP8EAjkAuQSBAGkEVgAyAzEAGQQRAC0E0QCWAfkAmwMPAF8EygCbBLgAjAH5AJsEEwAoA7AAUAO0ADwEygCbBM8AUAH5AJsC0gA8BJgAWgQ8ABkEiABuBF8AcwOxABkD1AAKBGYAlgQTACgFjgBkBSQAKAPyAJsD8gCbA/IAmwHjAFoDVgBaBoYAmwH5/6wEEwAoBBMAKAO0/1cDtP9XBEgALQWOAGQFjgBkBY4AZAWOAGQEgQBpBIEAaQSBAGkEVgAyAzEAGQQRAC0E0QCWAksAAANKAAAEuACMAksAAAQTACgDsABQA7QAPATPAFAC0gA8BJgAWgSIAG4EXwBzA9QACgRmAJYEEwAoBY4AZAUkACgB+QCbBFYAMgOwAFAEXwBzBJsAPAAA/9wAAP8lAAD/3AAA/lECjQCrAo0AoALaAEMDTQB5Aaj/ugAAAEYAAABGAAAARgAAAEYAAABIAAAARgAAAEYAAABGBDUBfAQ1AS4ENQC3BDUAgQQ1ASwENQC+BDUArwQ1AIEENQCaBDUA2wQ1AIUCjQDBBDUAswYAAQAGAAEAAkIANgYAAQAENQCeBDUAmAQ1AMsGAAEABgABAAYAAQAGAAEABgABAAAAAEYGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAUb/7oGAAEABgABAAYAAQAFtQA6BbUAOgH0/7oB9P+6BgABAAYAAQAGAAEABgABAASBADYENQA2BD3/ugQ9/7oD6QBKA+kASgZ/ABQHdgAUAyf/ugQe/7oGfwAUB3YAFAMn/7oEHv+6BRsAMgS1ACQDAP/3BgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEAAAAAMAAAAEYAAABGAAAAQAAAAEYGAAEABgABAAAA/9wAAP5RAAD/FgAA/xYAAP8WAAD/FgAA/xYAAP8WAAD/FgAA/xYAAP8WAAD/3AAA/xYAAP/cAAD/IAAA/9wEcwBKCAAAAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQACjQB/Ao0AXQYAAQAE7gAVA00AeQGoAA4B1v/cAagAVgHWABADdQAyA3UAMgGoAC0B1gATBRsAMgS1ACQB9P+6AfT/ugGoAJMB1gATBbUAOgW1ADoB9P+6AfT/ugJCAAADAP/3BbUAOgW1ADoB9P+6AfT/ugW1ADoFtQA6AfT/ugH0/7oEgQA2BDUANgQ9/7oEPf+6BIEANgQ1ADYEPf+6BD3/ugSBADYENQA2BD3/ugQ9/7oCswBfArMAXwKzAF8CswBfA+kASgPpAEoD6QBKA+kASgaSAD4GkgA+BD//ugQ//7oGkgA+BpIAPgQ//7oEP/+6CMkAPgjJAD4Gxf+6BsX/ugjJAD4IyQA+BsX/ugbF/7oEp/+6BKf/ugSn/7oEp/+6BKf/ugSn/7oEp/+6BKf/ugRaACoDmgA2BDX/ugMn/7oEWgAqA5oANgQ1/7oDJ/+6Bk8AJwZPACcCJP+6Ahr/ugSnAEYEpwBGAiT/ugIa/7oEzwAtBM8ALQMn/7oDJ/+6BA0ARwQNAEcBqP+6Aaj/ugK0ACMCtAAjAyf/ugMn/7oENQBFBDUARQH0/7oB9P+6AkIANgMA//cDmv+6Ayf/ugN1ADIDdQAyBRsAMgS1ACQFGwAyBLUAJAH0/7oB9P+6BFoAQATOAEkEWgAmBM4AOQRaAFMEzgBKBFoAUwTOAEoGAAEABgABAAAAAEYAAABGBgABAAYAAQAGAAEAAAAARgAAAEYGAAEABgABAAAAAEgAAABGBgABAAYAAQAGAAEAAAAARgAAAEYAAABGAAAARgAAAEAAAAAwBgABAAAAAEYAAABGBgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEAAo0AygKNAMcCjQDGBgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEAAQD/uggA/7oQAP+6BtwAYwU/AEQG1QChBVsAgwAA/dwAAPwvAAD8pgAA/lQAAPzXAAD9cwAA/ikAAP4NAAD9EQAA/GcAAP2dAAD79QAA/HIAAP7VAAD+1QAA/wIEGwCgBqwAawasABkAAP62AAD9cwAA/ggAAPymAAD+UwAA/REAAPvIAAD69AAA+q8AAPxyAAD7qgAA+2oAAPzxAAD8fQAA+90AAPzBAAD7mAAA/eoAAP6EAAD9wgAA/PEAAP1fAAD+dgAA/rwAAPzrAAD9bAAA/VgAAPyQAAD9FQAA/CwAAPwTAAD8EgAA+5YAAPuWAccAiAVW//0EcwBKBVb//QRzAEoFVv/9BHMASgVW//0EcwBKBVb//QRzAEoFVv/9BHMASgVW//0EcwBKBVb//QRzAEoFVv/9BHMASgVW//0EcwBKBVb//QRzAEoFVv/9BHMASgVWAKIEcwBLBVYAogRzAEsFVgCiBHMASwVWAKIEcwBLBVYAogRzAEsFVgCiBHMASwVWAKIEcwBLBVYAogRzAEsCOQBjAccAHwI5ALoBxwB8BjkAYwRzAEQGOQBjBHMARAY5AGMEcwBEBjkAYwRzAEQGOQBjBHMARAY5AGMEcwBEBjkAYwRzAEQG3ABjBT8ARAbcAGMFPwBEBtwAYwU/AEQG3ABjBT8ARAbcAGMFPwBEBccAoQRzAIMFxwChBHMAgwbVAKEFWwCDBtUAoQVbAIMG1QChBVsAgwbVAKEFWwCDBtUAoQVbAIMFVgAGBAAAIQVWAAYEAAAhBVYABgQAACEFVv/9BHMASgI5/+IBx/+wBjkAYwRzAEQFxwChBHMAgwXHAKEEcwCDBccAoQRzAIMFxwChBHMAgwXHAKEEcwCDAAD+/gAA/v4AAP7+AAD+/gRV//0C6wAMB2MABwVa//sEqQChA4AAhgSpAKEDgACGBccApARrAIgEc//9BAAAFARz//0EAAAUBVYACQQAAA8FVQBXBCsARQVVAKEEcwCHBgUAYwRzAFUGOQBgBHMARAW1ADoB9P+6AiT/ugIa/7oEpwBGAfQAngH0ABAB9AAbAfQAEAH0AGsB9P/5Aif/zgAAAA8AAP/1AqoApAKqAKQAAAAOAAAAVgAAAFYAAP/PAagADwHW/78BqP/1Adb/zQGoAB0B1v/1AagAkwHWABMDdQAyA3UAMgN1ADIDdQAyBRsAMgS1ACQFtQA6BbUAOgH0/7oB9P+6BbUAOgW1ADoB9P+6AfT/ugW1ADoFtQA6AfT/ugH0/7oFtQA6BbUAOgH0/7oB9P+6BbUAOgW1ADoB9P+6AfT/ugW1ADoFtQA6AfT/ugH0/7oFtQA6BbUAOgH0/7oB9P+6BIEANgQ1ADYEPf+6BD3/ugSBADYENQA2BD3/ugQ9/7oEgQA2BDUANgQ9/7oEPf+6BIEANgQ1ADYEPf+6BD3/ugSBADYENQA2BD3/ugQ9/7oEgQA2BDUANgQ9/7oEPf+6ArMAMgKzADICswBfArMAXwKzAF8CswBfArMAMgKzADICswBfArMAXwKzAF8CswBfArMAXwKzAF8CswA4ArMAOAKzAEkCswBJA+kASgPpAEoD6QBKA+kASgPpAEoD6QBKA+kASgPpAEoD6QBKA+kASgPpAEoD6QBKA+kASgPpAEoD6QBKA+kASgaSAD4GkgA+BD//ugQ//7oGkgA+BpIAPgQ//7oEP/+6BpIAPgaSAD4EP/+6BD//ugjJAD4IyQA+BsX/ugbF/7oIyQA+CMkAPgbF/7oGxf+6BKf/ugSn/7oEWgAqA5oANgQ1/7oDJ/+6Bk8AJwZPACcGTwAnAiT/ugIa/7oGTwAnBk8AJwIk/7oCGv+6Bk8AJwZPACcCJP+6Ahr/ugZPACcGTwAnAiT/ugIa/7oGTwAnBk8AJwIk/7oCGv+6BKcARgSnAEYEpwBGBKcARgk+ADIJPgAyB0D/ugdA/7oGfwAUB3YAFAMn/7oEHv+6BM8ALQTPAC0DJ/+6Ayf/ugTPAC0EzwAtAyf/ugMn/7oEzwAtBM8ALQMn/7oDJ/+6Bn8AFAd2ABQDJ/+6BB7/ugZ/ABQHdgAUAyf/ugQe/7oGfwAUB3YAFAMn/7oEHv+6Bn8AFAd2ABQDJ/+6BB7/ugZ/ABQHdgAUAyf/ugQe/7oEDQBHBA0ARwGo/7oBqP+6BA0ARwQNAEcBqP+6Aaj/ugQNAEcEDQBHAaj/ugGo/7oEDQBHBA0ARwGo/7oBqP+6BDUARQQ1AEUB9P+6AfT/ugQ1AEUENQBFBDUARQQ1AEUENQBFBDUARQH0/7oB9P+6BDUARQQ1AEUEgQA2BDUANgQ9/7oEPf+6AkIANgMA//cDGgAaAxoAGgMaABoDdQAyA3UAMgN1ADIDdQAyA3UAMgN1ADIDdQAyA3UAMgN1ADIDdQAyA3UAMgN1ADIDdQAyA3UAMgN1ADIDdQAyBRv/ugS1/7oFGwAyBLUAJAH0/7oB9P+6A3UAMgN1ADIFGwAyBLUAJAH0/7oB9P+6BRsAMgS1ACQGfwBFBn8ARQZ/AEUGfwBFAagAKAAA/ikAAP6iAAD/MAAA/x0AAP8SAAD/kgAA/n4I/AAyCK0AMgAA/7UAAP+2AAD+7QAA/2QAAP5+AAD/nwGNAAAC9v/9AAD+ggAA/xAEzQAyAAD/WAAA/1gAAP9kBpIAPgaSAD4EP/+6BD//ugjJAD4IyQA+BsX/ugbF/7oEWgAqA5oANgQ1/7oDJ/+6A00AeQK0ACMCQgA2AfT/ugKQ/7oB9AAvAfQAOwH0ABIB9ACxAfQAbQZ/ABQHdgAUAfkAmwAA/tkCvAAAA/IAmwRa//UEzv/1BFoAUwTOAEoEWgBTBM4ASgRaAFMEzgBKBFoAUwTOAEoEWgBTBM4ASgRaAFMEzgBKBDUAcQQ1AK0EWgAPBM4ADwRzABQGEQAUBUAApwRzAIYFQAAKBHMACgXHAFEFxwBmBAAAUAXH//0GegAUBUAASgRzAEYEdABIBVYAbgTVAFME4//EBjkAbQT+AA8HDACHAccAgwI5AB8FVgCWBAAAiAHHABUEAAAYByAApAXH/7gEcwCLBjkAYAbyAGMFVwBEBgkAFARzAIYFVgCeBVYAawQAAE8E8gCUAwsARAI5ACQE4wAUAjkAJATjADAF+wBhBccAoQYuABAEAAAhBOMAKQQAACgE4wApBOMAMQRcAEQEXAA/BHMAPARzAFUDqwAyA+UAJARzAIcCFAC8A04AvASsAHICOQCwCqoAngnHAJ4IZABGCH8AlgaqAJYDnACDCccAnAeOAJwGKwCHBHMAVQVW//0EcwBKAAD+/gVW//0EcwBKCAAAAQcdAEQGOQBtBHMAGgY5AG0EcwBCBVYAlgQAAIgGOQBjBHMARAY5AGMEcwBEBOMAKQRcAEwBx/+iCqoAngnHAJ4IZABGBjkAbQRzAEIIRgCkBPIAngXHAJwEcwCHBVb//QRzAEoFVv/9BHMASgVWAKIEcwBLBVYAogRzAEsCOf+KAjn/ZAI5AAQCOf/2BjkAYwRzAEQGOQBjBHMARAXHAKECqv/MBccAoQKqAGgFxwChBHMAdgXHAKEEcwCDBVYAXAQAAD8E4wAwAjkAJARcAFEDfgATBccApARzAIcFpgCkBNYAXgSGAF4E4wApBAAAKAVW//0EcwBKBVYAogRzAEsGOQBjBHMARAAA/v0GOQBjBHMARAY5AGMEcwBEBjkAYwRzAEQFVgAGBAAAIQRzAFcEcwBIBHMAhgRzAIYEAAATBAAAUARzAEYEcwBGBHMAVQXpAFUDqwBJA6sAMgUNADIEDwBEAjn/uQRzAEIEcwBCBHgAUAQCABkE7wAZBHMAiwRzAIcEcwCHAccAGQHHAFcC2QBEAp4AAAJuABQBxwCDBJMAgwaqAIQGqgCEBqoAhwRz/6YEcwCLBGwAhwRzAEQGUwBEBj8AVwRmAEQCqv/kAqr/5AKq/+QCqgCFAqoAhQKqAIUCqv/kBFUAigRVAIoEAAA/Acf/ogIU/7kBx/9yAssAAAI5AA8COQAkBHMAGQSMAFQEYACIBAAAGgXHAAYEAAAYBCgAGQQAACgEVAAoBFwATARcAHkEAAAkBAAAUAQAACQEAABQBjkAYwRAAIgEDwBJBHgAUARrAIgDLgAABAAACAM7AIgEcwBIBAAAJAQAAFAHtwBGB0AARggLAEYFswAkA28AJAXAACQGHAATBUoAgwUPAIMD4gAeBDgAYwMRAGQDEQBkAUb/zgHrAGQB6wAAAesAAALqAGQD2QAAApEAAAGHAFoC1wBeAccAgAHHAGwBxwCKAqoA+wKqAPsCygAyAsoAMgSsAHAErABwBKwAZQSsAGUCqgEhAqoA3gKqAFkCqgEhAqoAHQKqAFkCqgDeAjkAtgI5ALYCqgD7AqoA+wKqAKYCqgCmAqoApgKqAB0Cqv/iAqr/+wKUAAABQgBkArgAMgKgAAACygAyAxAAlgMQAJYDEACWAxAAlgMQAJYCqgBiAqoAYgKqACgCqgAdAqoARwRXAJYEVwCWBFcAlgRXAJYEVwBDBFcAQwRXAEMEVwBDBFcAQwMQAEMEVwAvBFcALwRXAC8EVwAvBFcALwMQAC8EVwAlBFcAJQRXACUEVwAlBFcAJQMQAC8EVwAaBFcAGgRXABoEVwAaBFcAGgMQABoEVwBCBFcAQgRXAEIEVwBCBFcAQgMQAEIEVwCWBFcAlgRXAJYEVwCWBFcAQgRXAEIEVwBCBFcAQgRXAEIDEABCBFcALwRXAC8EVwAvBFcALwRXAC8DEAAvBFcALwRXAC8EVwAvBFcALwRXAC8DEAAvBFcAJgRXACYEVwAmBFcAJgRXACYDEAAmBFcAQgRXAEIEVwBCBFcAQgRXAEIDEABCBFcAlgRXAJYEVwCWBFcAlgRXAEIEVwBCBFcAQgRXAEIEVwBCAxAAQgRXACYEVwAmBFcAJgRXACYEVwAmAxAAJgRXACMEVwAjBFcAIwRXACMEVwAjAxAAIwRXAC8EVwAvBFcALwRXAC8EVwAvAxAALwRXAEsEVwBLBFcASwRXAEsEVwBLAxAASwRXAJYEVwCWBFcAlgRXAJYEVwBCBFcAQgRXAEIEVwBCBFcAQgMQAEIEVwAaBFcAGgRXABoEVwAaBFcAGgMQABoEVwAkBFcAJARXACQEVwAkBFcAJAMQACQEVwAvBFcALwRXAC8EVwAvBFcALwMQAC8EVwBOBFcATgRXAE4EVwBOBFcATgMQAE4EVwCWBFcAlgRXAJYEVwCWAAD+wQAA/sYAAP2sAAD+2AAA/5IAAP7pAAD/TAAA/qAAAP7EAAD/zgAA/2YAAP6gAAD+2AAA/tgAAP+XAAD/mAAA/5kAAP/0AAD/QgAA/0IAAP9EAAD/XwAA/ocAAP/sAAD/pgAA/1EAAP9RAAD/UQAA/skAAP8cAAAAAAAA/ukAAP9MAAD/kwAA/yoAAP9WAAD/zgAA/ocAAP67AAD+xAAA/sQAAP7YAAD+2AAA/rMAAP7JAAD9rQAA/sgAAP6zAAD+yQAA/a0AAP4WAAD+5gAA/6YAAP6HAAD/RAAA/roAAP8jAAD/mgAA/awAAP6IAAAAAAAA/rAAAP+YAAD+kwAA/6YAAP6HAAD+HAAA/2YAAP9EAAD+sAAA/rAAAP6wAAD/AwAA/1IAAP0fAAD/UwAA/1MAAP9TAAD+tQAA/rUAAP/DAAD+rgAA/twAAP7HAAD+yAAA/twAAP4eAAD/QgAA/1EAAP63AAD+sAKqAN4CqgBZAqoA+gSaAHAEYAAABi4AFAeqAAAGLgAUBHsATAY/AFcEzwBEBjkAYwRzAEQFxwBwBAAAUATjAKgDOwCIBP8AAAQ8ADIGDQAKBJ0AQgcgAKQGqgCEBWUAYwRzAIsFZACkBAAACgVWAGsFVgBrBOAABQTFABkF5QBfBG4ARAO2ABQDRwAoBM8ARASVAFsEAABQAcf/ogY5AGADiQBNA4kAUAVWAKIFwAChBHMASwR4AIcKtABtBP4AEAY5ABQE5wAUB5kAvwW1AIgFWAABBAAABgcuAL8FkACIBqEAeAV7AHoIbQC/BvAAiATVAGYDqwAfBl8AOQWCAEgGOQBgBHMARAZtAAkFDAAaBm0ACQUMABoImABjBywARAaqACAE5gAcCYcAbQbQAFAAAP43CrQAbQT+ABAFxwBmBAAAUAQHABQAAP6mAAD+vAAA/5gAAP+YAAD8KwAA/EwFwAChBHgAhwVAAAQEKwAUBVYAngRzAIcFXQCkBGQAiATVAE4DqwAyBKkABAOAAAAF7wApBEkAKAcJAKQFLwCICRgAoAb2AIgGBgA+BCsAIwXHAGYEAABQBOMAMAOqACYHZwAxBYcAJgVVAFcEKwBFBuQACgVUAAoG5AAKBVQACgI5AL8HYwAHBVr/+wVXAKEEaACGBUAAEgSrABgFxwCkBGsAiAXHAKQEawCIBVUAVwQrAEUGqgCYBYAAjAKqAC4FVv/9BHMASgVW//0EcwBKCAAAAQcdAEQFVgCiBHMASwYFAGMEcwBVB2MABwVa//sE1QBOA6sAMgTVAE4EXABMBcAAoQR4AIcFwAChBHgAhwY5AGMEcwBEBjkAYARzAEQFwABKBBUAKwUVAAoEAAAhBRUACgQAACEFFQAKBAAAIQVVAFcEKwBFBxUAqAXAAIsFQABKBHMARge/AEoHAwBGB6YAZgaGAFMFTQBmBBMAUwfDABIHRwAYCEYApAcHAIgGOQBtBHgAUAX5ADAFUwAmAAD/QwAA/skAAP93AAD/sAAA/0cAAP9WAAD/dAAA/tcAAP6sAAAAAAAA/1IAAP9WAAAAAAAA/qwAAP2aAAAAAAAA/2oAAP98AAD/aQAA/1YAAP6sAAD/fwAA/1YAAP3vAAD/QwAA/2kAAP98AAAAAAAA/a4AAP+MAAABAgAA/v4AAP7+AAD+3wAA/t8AAP9YAAD/IAAA/v4FVv/9BHMASgVWAJYEcwCGBVYAlgRzAIYFVgCWBHMAhgXHAGYEAABQBccAngRzAEYFxwCeBHMARgXHAJ4EcwBGBccAngRzAEYFxwCeBHMARgVWAKIEcwBLBVYAogRzAEsFVgCiBHMASwVWAKIEcwBLBVYAogRzAEsE4wCoAjkAEwY5AG0EcwBCBccApARzAIcFxwCkBHMAhwXHAKQEcwCHBccAkwRzAGgFxwCkBHMAhwI5/98Bx/+SAjkAIAI5AAYFVgCWBAAAiAVWAJYEAACIBVYAlgQAAIgEcwCWAccAfgRzAJYBx/+5BHMAlgHH/6UEcwCWAcf/owaqAJgGqgCHBqoAmAaqAIcGqgCYBqoAhwXHAJwEcwCHBccAnARzAIcFxwCcBHMAhwXHAJwEcwCHBjkAYwRzAEQGOQBjBHMARAY5AGMEcwBEBjkAYwRzAEQFVgCeBHMAhwVWAJ4EcwCHBccAoQKqAIUFxwChAqoAhQXHAKECqgBeBccAoQKqACYFVgBcBAAAPwVWAFwEAAA/BVYAXAQAAD8FVgBcBAAAPwVWAFwEAAA/BOMAMAI5ACQE4wAwAjkAJATjADACOf//BOMAMAI5AA4FxwChBHMAgwXHAKEEcwCDBccAoQRzAIMFxwChBHMAgwXHAKEEcwCDBVYACQQAABoFVgAJBAAAGgeNABkFxwAGB40AGQXHAAYFVgAJBAAADwVWAAkEAAAPBVYABgQAACEE4wApBAAAKATjACkEAAAoBOMAKQQAACgEcwCHAjkAAwXHAAYEAAAhBHMASgHHAIkEoABIBKAASASgAEgEoABIBKAASASgAEgEoABIBKAASAVW//0FVv/9BoIAEwaCABMGggATBoIAEwaCAFYGggBWA5EAYgORAGIDkQBiA5EAYgORAGIDkQBiBh4AAAYeAAAHbAAAB2wAAAdsAAAHbAAABHMAiwRzAIsEcwCLBHMAiwRzAIsEcwCLBHMAiwRzAIsGjwAABo8AAAgfAAAIHwAACB8AAAgfAAAIH//zCB//8wHHAIEBxwCBAcf/mwHH/5sBx//rAcf/6wHH/6IBx/+iAwEAAAMBAAAEkQAABJEAAASRAAAEkQAABJH/8wSR//MEcwBEBHMARARzAEQEcwBEBHMARARzAEQGnQAABp0AAAgtAAAILQAAB8kAAAfJAAAEYACIBGAAiARgAIgEYACIBGAAiARgAIgEYACIBGAAiAaCAAAHrgAACBIAAAeuAAYGPwBXBj8AVwY/AFcGPwBXBj8AVwY/AFcGPwBXBj8AVwZfAAAGXwAAB+8AAAfvAAAHiwAAB4sAAAeL//8Hi///BKAASASgAEgDkQBiA5EAYgRzAIsEcwCLAcf/5gHHAGgEcwBEBHMARARgAIgEYACIBj8AVwY/AFcEoABIBKAASASgAEgEoABIBKAASASgAEgEoABIBKAASAVW//0FVv/9BoIAEwaCABMGggATBoIAEwaCAFYGggBWBHMAiwRzAIsEcwCLBHMAiwRzAIsEcwCLBHMAiwRzAIsGjwAABo8AAAgfAAAIHwAACB8AAAgfAAAIH//zCB//8wY/AFcGPwBXBj8AVwY/AFcGPwBXBj8AVwY/AFcGPwBXBl8AAAZfAAAH7wAAB+8AAAeLAAAHiwAAB4v//weL//8EoABIBKAASASgAEgEoABIBKAASASgAEgEoABIBVb//QVW//0FVv/9BVb//QVW//0CqgDlAqoA/QKqAOUCqgAGAqoABgRzAIsEcwCLBHMAiwRzAIsEcwCLBoIAAAaCAAAG8wAABvMAAAXHAKQCqgATAqoAEwKqAAYBx/+7Acf/qwHH/8oBx//KAcf/kwHH/5MCOQAaAjn/9QNlAAADZQAAAqoAEwKqABMCqgAGBGAAiARgAIgEYACIBGAAiASNAIMEjQCDBGAAiARgAIgFVgAGBVYABgbmAAAHGAAABh4AAAKq/+oCqv/qAqoAWQY/AFcGPwBXBj8AVwY/AFcGPwBXB2UAAAadAAAHJwAABl8AAAX7AGECqgDeAqoA5QRzAA0FxwBmBccAZgaqAIcFxwAkCVAAoQeNABkFVgAfBOMAMAgAACkEAAAwBMEAZgAA/1MAAP9TAAD/UwAA/1MBxwAZAcf/ogQrAAUFVgARBXQARgLL/6MFegCHAvD/yAV/AAoFfwAKAqoAhAKqAIQCqgDJAqoAyQKqAKACqgBZAqr/rwKqADoCqgAGAjkAuQKqAKkCqgCpAqoAqQKqAKkDLgAeAy4AHgKqADoAAP9zAAD/pQAA/tgAAP8jAAD/cgAA/3IAAP7nAAD/pQAA/1MAAP9TAAD/UwVWAJ4EcwCHA/gAGQX7ABkHHQBEBEAAGQQAAFAEaQCHBGkAGQPrAIcDqwAyAccAiANhAEEEAACIAzYAEAWAAIwEeACHBHMARAQAABME3gBEBN4ARATeAA0HjQBQA6gARARzAEQEcwBEBCsAhARVAB8EVQAfA6oAJgRgAIgExgBEBd4ARATGAEQEAAAaBccABgQAACgDqwAyA2sAPwTbAB8C6wCIBAAAGgRVAIgEKwCEBbQAegSrABgDoAAABU8AAANRADIDUf/RA5gAMgNIADIDSAAyA/gAMgNuADIBVgBpAoQALQNmADIC0AAyBBUAMgNxADIDbwAyBBgAMgMPADIDWQAyA5wAMgN2ADEDbwAyBPsAAAL6ADIC+gAyAwQAMgTMADIDBQBkAwUAMgL5ADIC+QAyAowAMgKMADIDBAAyAUIAZAK2AGQElQBkAw8AZAMFADIC1QAyAwUAMgMFADIDBgBkAcIAMgMPAGQDQgAyBJUAZAKSAAADIAAAAxUAZAKSAAADBgAyA4UAMgK/AAABQgBkAesAZAMPAGQCkgAAAxUAZAKSAAADCQAyA4UAMgK/AAAF7QBGCmYARgYTAEYGif+6BUH/ugHpADwEWgARAAD/DQAA/zUAAP7OAAD+twAA/skAAP/PAAD/TwAA/54AAP7KArMAXwKzAF8D6QBKA+kASgOa/7oDJ/+6A5r/ugMn/7oFrQBpBT0ALQX9AJYE3ABQBOAAPAX2AJsFPwAoBlAAKASsAHIAAP47AAD+ZgAA/mYEc//8AqoAUwLV/84BqP+6Aaj/ugGo/7oBqP+6BlgAFQnFAEcEAAAACAAAAAQAAAAIAAAAAqsAAAIAAAABVQAABHMAAAI5AAABmgAAAKsAAAAAAAAF5QADBccAZgaqAJgFgACMB0QAgwcYAEYHGABIBVb//QXHAGYEAAAUBHMACgTjADAEAABPBAAAKASlAB0AAAECAAD/QgAA/r8AAP86AAD/UwSNAAoFxwBRBccAZgXHAFEEVQChAusAiAAA/0MAAP8EAAD/rALSAJYAAP83Ahr/ugJQAB4AAP86AAD/WwAA/18AAP9+AAD/lAAA/0oAAP6cBbUAOgW1ADoB9P+WAfT/lgW1ADoFtQA6AfT/ugH0/7oFtQA6BbUAOgH0/7oB9P+6BbUAOgW1ADoB9P+6AfT/ugW1ADoFtQA6AfT/ugH0/7oFtQA6BbUAOgH0/7oB9P+6BbUAOgW1ADoB9P+6AfT/ugSBADYENQA2BD3/ugQ9/7oEgQA2BDUANgQ9/7oEPf+6ArMAMgKzADICswBfArMAXwPpAEoD6QBKBpIAPgaSAD4EP/+6BD//ugRaACoDmgA2BDX/ugMn/7oEWgAqA5oANgQ1/7oDJ/+6BFoAKgOaADYENf+6Ayf/ugZPACcGTwAnAiT/ugIa/7oGTwAnBk8AJwIk/7oCGv+6Bn8AFAd2ABQDJ/+6BB7/ugZ/ABQHdgAUAyf/ugQe/7oGfwAUB3YAFAMn/7oEHv+6ArQAIwK0ACMDJ/+6Ayf/ugK0ACMCtAAjAyf/ugMn/7oENQBFBDUARQH0/7oB9P+6BDUARQQ1AEUB9P+6AfT/ugQ1AEUENQBFAfT/ugH0/7oEDQBHBA0ARwGo/7oBqP+6A+kASgPpAEoD6QBKA+kASgaSAD4GkgA+BD//ugQ//7oEc/+TBHMARgI5/78Gqv/VBHP/twRz/5ECqv+kAqr/pAQA//8COf+5BAAAKARzAIkDCwBkBHQASAZJACQBxwAZAccAGQRzAB4EYAAeBIwACgRzAIYEcwBGAjkAEwW0AEIEAACIAcf//AaqAIcEcwCLBHMAhwKq//sEAAA/Axj/ogQAABoEAAAPBAAAKARzAEoEcwBIBHMARgRzAEsDqwBJA6sAMgU0AFUBxwCIBAAAEwHH/6IEcwCDBFwATAMEAGQC1QAyAskAMwL8ADICjAAyAdUAMgHVAAADBAAyAxEAZAFCABkBQgBkAUIAZAFCABkCKgAAAUIAZAFCAAkCMwBkBJMAZASTAGQDD//JAw8AZAMOAGQDBQAyAwAAMgK4ADIBQv/KAcIAMgMPAB0DGgAyAwYAZALUAGQCkgAAAt4AMgLeADIC3gAyAvQAMgLqADIAAP68AAD+vAAA/3MAAP6pAjkAuQL6ADIC+QAyAwUAMgKgAAAC+QAyBjkAbQVW//0EcwAPBccAZgKqAEEEoABIBKAASASgAEgEoABIBKAASASgAEgEoABIBKAASAHH/5sBx/+rAcf/mwHH/6sBx/+bAcf/uwHH/5sBx/+7BGAAiARgAIgEYACIBGAAiARgAIgEYACIBGAAiARgAIgBx/+rAcf/qwHH/7sBx/+7BGAAiARgAIgEYACIBGAAiARaAFMEzgBKA6AAEwVWABEFxwApBVgACwVWAKIEcwBLBAAAMwHH/6IF5gBjBHMASAXHAAACqgAPBVYABgQAACEEAAATBAAAUAQAABMBxwCDBFX//QLrAAEFVgAJBAAADwVWAAkEAAAPBNUAUwOrAEkFQAASBKsAGAAA/sYAAP7UAAD+xgAA/tQAAP5fAAD+XwAA/3IAAP9zAAD+5weLAAoD6wBMBAAAEwRzAAoBxwAVBHP/9AVWABEFxwChBHMAGQI5/4sFxwCkBHMAhwVWAJYEAACIBOMAKQQAACgEAAA7BJ4ApANnAIgFMABIAAD/UwAA/7wAAP7+AAD+/gAA/qQAAP6kAccAiAXJAKUFxwCcBckApQAA/s0AAP9IAAD+yQAA/s4AAP7FAAD+0AAA/tEAAP7uAAD+1gAA/twAAP3ZBjkAWARzAEgHjQAZBccABgWfAKQAAP65BdwAYwTGAAkITAAZBroABgI5ALkDgAByAYcAWgGHAFoEAACZBAAAmQI5ALACOQCwAjkAsAKqABkE4wAwBHMAUARzAA8EcwAcBlsAhwZKAEwAAAAAAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAHSAAAB0gAAAdIAAAJSAAAC+AAAAvgAAANgAAAD2AAABB4AAARaAAAEygAABoYAAAdiAAAJjAAAC2YAAAzGAAAOgAAAEFYAABECAAATlgAAFcoAABYmAAAWJgAAFiYAABaWAAAWlgAAF4gAABeIAAAZMgAAGsoAABwEAAAdTAAAHhAAAB7GAAAgVgAAIVwAACJAAAAiQAAAIkAAACLKAAAl9AAAJ54AACjSAAAp2AAAK8wAAC44AAAw4gAAMZAAADK0AAA0KAAANmYAADlyAAA7GAAAPFgAADxYAAA8WAAAPFgAADxYAAA8jAAAPIwAAD9eAABBPAAAQvAAAESkAABGYgAAR7YAAEmmAABLSgAATD4AAEw+AABO1gAAT9IAAFICAABTyAAAVYoAAFdOAABY5AAAWeoAAF2SAABetgAAYFQAAGJyAABm3AAAaQAAAGtYAABtQAAAbUAAAG1AAABtQAAAbUAAAG1AAABtQAAAbUAAAG1AAABtQAAAbUAAAG1AAABtQAAAbUAAAG1AAABtQAAAbUAAAG1AAABtQAAAbUAAAG1AAABtQAAAbUAAAG1AAABtQAAAbUAAAG1AAABtQAAAbUAAAG1AAABtQAAAbUAAAG1AAABtQAAAbUAAAG1AAABtQAAAbUAAAG1AAABtQAAAbUAAAG1AAABtQAAAbUAAAG1AAABtQAAAbzAAAG8wAABvMAAAbzAAAG8wAABvMAAAbzAAAG8wAABvMAAAbzAAAG8wAABvMAAAbzAAAG8wAABvMAAAbzAAAG8wAABvMAAAbzAAAG8wAABvMAAAbzAAAG8wAABvMAAAbzAAAG8wAABvMAAAbzAAAG8wAABvMAAAbzAAAG8wAABvMAAAbzAAAG8wAABvMAAAbzAAAG8wAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAAAb2gAAG9oAABvaAABAAANXQDyADwAnQAHAAIAEAAvAFYAAASs//8ABQACAAAAFAD2AAEAAAAAAAAAEAAAAAEAAAAAAAEADAAQAAEAAAAAAAIABwAcAAEAAAAAAAMADAAjAAEAAAAAAAQADAAvAAEAAAAAAAUADAA7AAEAAAAAAAYADABHAAEAAAAAAAcABwBTAAEAAAAAAAgABwBaAAEAAAAAAAkABwBhAAMAAQQJAAAAIABoAAMAAQQJAAEAGACIAAMAAQQJAAIADgCgAAMAAQQJAAMAGACuAAMAAQQJAAQAGADGAAMAAQQJAAUAGADeAAMAAQQJAAYAGAD2AAMAAQQJAAcADgEOAAMAAQQJAAgADgEcAAMAAQQJAAkADgEqT3JpZ2luYWwgbGljZW5jZUJPR0FJQStBcmlhbFVua25vd25CT0dBSUErQXJpYWxCT0dBSUErQXJpYWxWZXJzaW9uIDAuMTFCT0dBSUErQXJpYWxVbmtub3duVW5rbm93blVua25vd24ATwByAGkAZwBpAG4AYQBsACAAbABpAGMAZQBuAGMAZQBCAE8ARwBBAEkAQQArAEEAcgBpAGEAbABSAGUAZwB1AGwAYQByAEIATwBHAEEASQBBACsAQQByAGkAYQBsAEIATwBHAEEASQBBACsAQQByAGkAYQBsAFYAZQByAHMAaQBvAG4AIAAwAC4AMQAxAEIATwBHAEEASQBBACsAQQByAGkAYQBsAFUAbgBrAG4AbwB3AG4AVQBuAGsAbgBvAHcAbgBVAG4AawBuAG8AdwBuAAAAAwAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAALkAVAMosyYYH9C8AykA4AMpAAIDKbIrHR+5AycDHbI7H0C4AyOzEhUyD0EtAyAAAQAvAyAAAQAgAyAAbwMgAK8DIAC/AyAABABfAx4AAQAQAx4AfwMeAIADHgCvAx4AvwMeANADHgAGAAADHgAQAx4AIAMeAG8DHgCfAx4A4AMeAAYDHQMcsiAfEEEnAxkAfwMZAAIADwMXAO8DFwD/AxcAAwAfAxcALwMXAE8DFwBfAxcAjwMXAJ8DFwAGAA8DFwBfAxcAbwMXAH8DFwC/AxcA8AMXAAYAQAMXspIzQLgDF7KLM0C4AxezamwyQLgDF7JhM0C4AxezXF0yQLgDF7NXWTJAuAMXs01RMkC4AxezREkyQLgDF7I6M0C4AxezMTQyQLgDF7MuQjJAuAMXsycsMkC4AxezEiUygLgDF7MKDTLAQRYDFgDQAxYAAgBwAxYAAQLEAA8BAQAfAKADFQCwAxUAAgMGAA8BAQAfAEADErMkJjKfvwMEAAEDAgMBAGQAH//AAwGyDREyQQoC/wLvABIAHwLuAu0AZAAf/8AC7bMOETKfQUoC4gCvAuIAvwLiAAMC4gLiAuEC4QB/AuAAAQAQAuAAPwLgAJ8C4AC/AuAAzwLgAO8C4AAGAuAC4ALfAt8C3gLeAA8C3QAvAt0APwLdAF8C3QCfAt0AvwLdAO8C3QAHAt0C3QAQAtwAAQAAAtwAAQAQAtwAPwLcAAIC3ALcABAC2wABAtsC2wAPAtoAAQLaAtr/wALTsjc5Mrn/wALTsisvMrn/wALTsh8lMrn/wALTshcbMrn/wALTshIWMrgC0rL5KR+5AyYDHLI7H0C7AyIAPgAzAyKyJTEfuAMYsjxpH7gC47MgKx+gQTAC1ACwAtQAAgAAAtQAEALUACAC1ABQAtQAYALUAHAC1AAGAGAC1gBwAtYAgALWAJAC1gCgAtYAsALWAAYAAALWABAC1gAgAsoAIALMACAC1gAwAtYAQALWAFAC1gAIAtCyICsfuALPsiZCH0EWAs4CxwAXAB8CzQLIABcAHwLMAsYAFwAfAssCxQAXAB8CyQLFAB4AHwLKAsayHh8AQQsCxgAAAscAEALGABACxwAvAsUABQLBsyQSH/9BEQK/AAEAHwK/AC8CvwA/Ar8ATwK/AF8CvwCPAr8ABgK/AiKyZB8SQQsCuwDKCAAAHwKyAOkIAAAfAqYAoggAQGofQCZDSTJAIENJMkAmOj0yQCA6PTKfIJ8mAkAmlpkyQCCWmTJAJo6SMkAgjpIyQCaEjDJAIISMMkAmeoEyQCB6gTJAJmx2MkAgbHYyQCZkajJAIGRqMkAmWl8yQCBaXzJAJk9UMkAgT1QyuAKetyQnHzdPawEgQQ8CdwAwAncAQAJ3AFACdwAEAncCdwJ3APkEAAAfApuyKiofuAKaQCspKh+AugGAvAGAUgGAogGAZQGAfgGAgQGAPAGAXgGAKwGAHAGAHgGAQAGAuwE4AAEAgAFAtAGAQAGAuwE4AAEAgAE5QBgBgMoBgK0BgHMBgCYBgCUBgCQBgCABN0C4AiGySTNAuAIhskUzQLgCIbNBQjJAuAIhsz0+Mg9BDwIhAD8CIQB/AiEAAwC/AiEAzwIhAP8CIQADAEACIbMgIjJAuAIhsxkeMkC4AiKzKj8yQLgCIbMuOjJvQUgCwwB/AsMAjwLDAN8CwwAEAC8CwwBgAsMAzwLDAAMADwLDAD8CwwBfAsMAwALDAO8CwwD/AsMABgDfAiIAAQCPAiIAAQAPAiIALwIiAD8CIgBfAiIAfwIiAO8CIgAGAL8CIQDvAiEAAgBvAiEAfwIhAK8CIQADAC8CIQA/AiEATwIhAAMCwwLDAiICIgIhAiFAHRAcECsQSAOPHAEPHgFPHv8eAjcAFhYAAAASEQgRuAENtvcN+PcNAAlBCQKOAo8AHQAfApACjwAdAB8Cj7L5HR+4AZiyJrsfQRUBlwAeBAEAHwE5ACYBJQAfATgAcwQBAB8BNQAcCAEAHwE0ABwCqwAfATKyHFYfuAEPsiYsH7oBDgAeBAG2H/kc5B/pHLgCAbYf6By7H9cguAQBsh/VHLgCq7Yf1ByJH8kvuAgBsh+8JrgBAbIfuiC4AgG2H7kcOB+tyrgEAbIfgSa4AZqyH34muAGath99HEcfaxy4BAGyH2UmuAGash9ec7gEAUAPH1ImWh9IHIkfRBxiH0BzuAgBth8/HF4fPCa4AZqyHzUcuAQBth8wHLsfKxy4BAG2HyocVh8pHLgBAbIfIx64BAGyH1U3uAFoQCwHlgdYB08HNgcyBywHIQcfBx0HGwcUCBIIEAgOCAwICggICAYIBAgCCAAIFLj/4EArAAABABQGEAAAAQAGBAAAAQAEEAAAAQAQAgAAAQACAAAAAQAAAgEIAgBKALATA0sCS1NCAUuwwGMAS2IgsPZTI7gBClFasAUjQgGwEksAS1RCsDgrS7gH/1KwNytLsAdQW1ixAQGOWbA4K7ACiLgBAFRYuAH/sQEBjoUbsBJDWLkAAQERhY0buQABASiFjVlZABgWdj8YPxI+ETlGRD4ROUZEPhE5RkQ+ETlGRD4ROUZgRD4ROUZgRCsrKysrKysrKysrGCsrKysrKysrKysrGCsdsJZLU1iwqh1ZsDJLU1iw/x1ZS7CTUyBcWLkB8gHwRUS5AfEB8EVEWVi5Az4B8kVSWLkB8gM+RFlZS7gBVlMgXFi5ACAB8UVEuQAmAfFFRFlYuQgeACBFUli5ACAIHkRZWUu4AZpTIFxYuQAlAfJFRLkAJAHyRURZWLkJCQAlRVJYuQAlCQlEWVlLuAQBUyBcWLFzJEVEsSQkRURZWLkXIABzRVJYuQBzFyBEWVlLuAQBUyBcWLHKJUVEsSUlRURZWLkWgADKRVJYuQDKFoBEWVlLsD5TIFxYsRwcRUSxHhxFRFlYuQEaABxFUli5ABwBGkRZWUuwVlMgXFixHBxFRLEvHEVEWVi5AYkAHEVSWLkAHAGJRFlZS7gDAVMgXFixHBxFRLEcHEVEWVi5DeAAHEVSWLkAHA3gRFlZKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKytlQisrAbM7WWNcRWUjRWAjRWVgI0VgsIt2aBiwgGIgILFjWUVlI0UgsAMmYGJjaCCwAyZhZbBZI2VEsGMjRCCxO1xFZSNFILADJmBiY2ggsAMmYWWwXCNlRLA7I0SxAFxFVFixXEBlRLI7QDtFI2FEWbNHUDQ3RWUjRWAjRWVgI0VgsIl2aBiwgGIgILE0UEVlI0UgsAMmYGJjaCCwAyZhZbBQI2VEsDQjRCCxRzdFZSNFILADJmBiY2ggsAMmYWWwNyNlRLBHI0SxADdFVFixN0BlRLJHQEdFI2FEWQBLU0IBS1BYsQgAQllDXFixCABCWbMCCwoSQ1hgGyFZQhYQcD6wEkNYuTshGH4bugQAAagACytZsAwjQrANI0KwEkNYuS1BLUEbugQABAAACytZsA4jQrAPI0KwEkNYuRh+OyEbugGoBAAACytZsBAjQrARI0IAK3R1c3UAGEVpREVpREVpRHNzc3N0dXN0dSsrKyt0dSsrKysrc3Nzc3Nzc3Nzc3Nzc3Nzc3Nzc3Nzc3NzcysrK0WwQGFEc3QAAEuwKlNLsD9RWlixBwdFsEBgRFkAS7A6U0uwP1FaWLELC0W4/8BgRFkAS7AuU0uwOlFaWLEDA0WwQGBEWQBLsC5TS7A8UVpYsQkJRbj/wGBEWSsrKysrKysrKysrKysrKysrK3UrKysrKysrQ1xYuQCAAruzAUAeAXQAc1kDsB5LVAKwEktUWrASQ1xaWLoAnwIiAAEAc1kAK3RzASsBcysrKysrKysrc3NzcysrKysrACsrKysrKwBFaURzRWlEc0VpRHN0dUVpRHNFaURFaURFaURzdEVpREVpRHMrKysrK3MrACtzK3R1KysrKysrKysrKysrKytzdHVzK3N0dXN0dSsrK3QrKwAA); }&#xA;@font-face { font-family: &quot;g_font_6&quot;; src: url(data:font/opentype;base64,T1RUTwAJAIAAAwAQQ0ZGINnUzR0AAACcAAAYDE9TLzJEqqxTAAAYqAAAAGBjbWFwIZficwAAGQgAAAB8aGVhZKsnT+UAABmEAAAANmhoZWED8QHJAAAZvAAAACRobXR4A/cAAAAAGeAAAAEMbWF4cABDUAAAABrsAAAABm5hbWVPS2/FAAAa9AAAAgpwb3N0AAMAAAAAHQAAAAAgAQAEAgABAQEPQk9HQkREK0FyaWFsTVQAAQEBJv0t+9kcB9D6ggUdAAAAUA8dAAAAbxEdAAAACR0AABgCEvgbDBYAAQEBCEFyaWFsTVQAAAABAAEAAAkBAAwAAA8AABEJACIIACwPAEIIAEwPAG8AAEMCAAEAGAAbAFsAnAC3AMEBSgFyAewCoALFAzgD7gQhBPgFtwXtBqAHKwejB7wH0gh2CI8ImwjGCNMJCwkoCbAKDQq4C0AMGQwrDIEMqg0EDU8NgA2kDn8O8A9mD+AQXBCeEUkRlBGqEdQR4BJkErQTIxOmFBsUWBUkFXMVyhX0FjAWbRbTFv4XCcb5BRb5BfyI/QUHm/j1Ffho/OX8aAYO/DEO+/r3vftmFSr3MFr3MfcwGsiSyZnIHpa7m7qfuJiopbuyzwhMBk45XjluOQhyRH5BPRo0nDasOR6tObRDu04IDvv694uQFazdnODiGtl+1XLSHm7dXt1O3QhMBrNHpVqYbp5em1yWWgiZT5JOThr7MFr7MSr7MB7KBrvItNOt3QgOIPfi9wgV91j3V937V/dXOPtX+1c591f7WAcO/DH3UxbvJycHDvcFyRVassFy0Bu/t5mnrR+tp6WznL8InL6Uz98a0obEgLQegLV8r3moeKhzoW6bCJpuaZNlG1dgfW9pH2hvcWR6Vwh6V4JHNhr7GqMquk8ey/ipFa2jrJyzG7SteGSnH6ZkmT37Chr7Cn09cGQeZG9peGMbY2mesm8fcLJ92fcKGvcKmtuptx4O+Aj5YxVSBnxscWtmamZqYG9adAg2B6aVqpuun62fp5+gnwj8xOMHDvcr3xWVm5ibmpuamq2qv7fLwLi1pqqmqp+olqYIl6eRp6gaw3e7Y7EesWNUnkcbR1R5aGMfYmh0V4VI5YIYuJiupaQepKStmLYbs6x/c6QfpHOXbmgaan1ncGYeb2ZWWD5LWWNlZ3BrcGx4a35rhHiHdox2CPhu3wYO9wW3FWa1v3jKG9DFoba5H7i3osDJGrp/sXSqHnSqap9glayao5+cpAicpJOoqRqsgqp6px55qHKiapwInGpok2MbU1t7amUfZWtzXYBQ43sYkraZrKKhCKCip5auG62ngHahH6F2lnFqGmN8bW13HnhtaYFmG4eGi4yFH4I+BZKjoI6cG7OtfnClH6ZxmGpjGmB9aG5uHm5vaH1hG2htlqFzH3Oheq+BvTN/GJFPo1u0ZQgO+C8W9z/s3Cr4ZEMH+9v8ZAU698v7Pwf7dfeQFfd199YF+9YHDvcEthVmtcB5zBvayqjFuB+xup7DzBrPdsNgth62YFahTRtcXnxtYB+x91UF97Hf+/cGRvwE3n+YoJ2coZgZmKKkkagbubB9bqYfp26ZY1kaVnxhbmsea25ne2EbZ22WonIfc6F7rYS4L4QYkU+iWrRnCA74Rvk0FapnXZtSG0BPcFReH1hMcSf7Hxr7EKIzuVUeVbrGcNUbtrGVoK0frZ+mqZ6xCJ6ylbW4Gs92w2K2HrZiWaFQG2pqg3xtH2x7cXN2a4zSk8ObsZuyoaimoAiaoaSTpxuuqX5yox+ZfJZyk2jikhiEw3W2Z6sI+5H73BWopq2ZsxuzrH1uph+lb5hkWRpYfmJwbR5tcWt8ZRtxc5KadB90mXmgfqcIfqeFqKkauZmxp6ceDvgh+QMVXlhhTWRAZEFsPnY7djyARopTCOUGkNKWzZ3Ho+Cu3rfbuNy4zLm7CM/8YzcHDtf32BV0bH9kXBpNoVe2YR5htsR20hvRxKC0th+2taG/yBq3gLF0qx50q2qiX5mumaaenKMInKSUqKwav3i3ZbAer2VZnUwbTVl5aGYfZmd4X1caaZRtnHIenXOmeLB9X4BpdXNsCPcJ97cVoKGnlq0brKeAdaEfoXWWcGsabIBwdnYednVwgGgbaG+WoHUfdqGAp6waqZaloaEedfvGFaamrpm0G7aufXCnH6dvmWhhGmF9aXBwHnBwaH1hG3BykZhzH3SYeZ2Aowh/ooWjpBq0mK6mph4O9wuuFWyuuXvDG8C5maeyH7KoqLSfwQifwZXU5xrjgc53uR53um6uZKQIpGVgmF0bSlZ1X2AfYF52UUIaRZ9StGAeYLS9dsYbr6yUnKkfqp2ioZ2nCIOMhocaZoZngmgeg2iAb352fnd6end/CH52dIVwG2txlJ13H3edfaeEszeEGJJToF+vbAj3lPfdFW5xaX1jG2JpmahwH3CnfbC4Gr6ZtKirHquorZuyG7GrfG6mH6ZtmGNZGlh+ZHFvHg5z7hbZ920F98EG3vttBfcABvu4+WAFIwb7p/1gBfex+IwVm7iZuZW6lmScWaJO1vtaGPuIBg5z9+4WubGPk6sfqpOll6CaoJudoZmoCJmokqqtGrR/r3SqHnSqaaBgmK2cpKCbpgicppOoqhqsgqp4qR54qXGiapkImmpfklUb+6H9YAbq+QwV9yMGv6+IhKAfoIScf5Z5CJZ5kXZzGnKFdn96Hn56eYBzgwiGeW2IYRv7LwY3BPc6Briuh4OjH6SDnn2YdwiZeJJzcRp0hnaCeh6BeX9+fYJ8gnmEdYcIiX91imwb+0YGDqr4lfcHFWxmXnxWG2BilqJmH2ahb616uAh5uYLAyBq6krmatx6auKWusKUIprC5mMIbu7J/c6sfqnSjZZxX6KEYeM1pvlqvCLBaT51EG0tSfW5WH1duYmFvUwhuVH1KQBpHmEukUB6kT7Beu2sIbLvKe9gb1cqftL8fvrSvxp/ZLKMYfk9yXWdtCA6q9+MWt7GPk6wfrZOnl6Obo5ugoZ+mn6ebrZi1CJi1kbzBGsuCw3i9Hni9b7Rlqm6kaJxilQiSbmCOVBv7i/1gBur5DBX3KgbDtIaBpR+ufqlwo2IIpGOXUUAaVYVdfmUef2V5bXV0e3t1f3GCCIJwZodcG/stBg5z+PkW3/xL94j4H9/8H/dw+Drf/Jn9YAcOO/dFFvfZ9+Tf++T3c/gY3/x3/WAHDuL5AvetFfsaB3d5bXpkewh7ZGODYhtcX5WgYR9hoGurdbYIdbaAwcsav5S7nbcelqWao56gn6GknKuYCJiqsZK2G6+shX6oH6l/onqbdpt2mG+WZuCjGH+7ebJzqXOpaqJinAicYVyTVxtETHxuVB9VbmFebk8Ibk58SkYaRJpMqFIeqFK3X8RtCG3Ey3zSG7++lJ68H7yeu6e6sAj3nfvDNwcOqvdEFvfl+Ab75er5YCz7u/wG97ss/WAHDvwx91AW+WAs/WAHDnP3PBb3jAf3CfcF95P7/QX3EQb7zfg+98D3tgX7FAb7+Pv3Bff3LP1gBw74nBbf+/T5DCz9YAcO9yL3Ohb49gf3Y/z2BeAG92X46wX86+b5YPsTB/tA/IZ5WH9lg3EZg6OArnu6+z34jxj7Iv1gBg6q9zsW+MYH+Az8xgXs+WAw/MYG/Az4xgUq/WAGDuLk9z4VplO0XsBrCGrAx3vPG8nFmqjAH8GptbaoxAioxJrM1BrSfctvxB5vw2O3VqsIqlZPm0kbJjlpSEsfS0hrLvsLGk2ZT6ZTHvcV+CsVubzEos4bu7V/c7EfsXOoap5fCJ9glVhRGi90RF1ZHlldUHJEG0VRpLxdH1y9dM/hGvaj2Lu5Hg5z90AW97j3TAfw0aC1sh+ytZ6/xxqvhKt8qR59qHiic5xzm26WZ5EIkHJnjVsb+6L9YAbq+QwV90sGtqmJh5ofpISffZp1CJp2k3FtGmJ+a3F0HnRyX4BOG/tNBg7i+VD3WxWdupTAxhrSfctvwx5vxGO3VqoIqlZQm0gbSlB8bVYfVmxjX25RCG5SfUpFGkSZS6hTHqdStF+/bAhswMZ7yxvLxpqowB++Y75uv3mnzBhmmWKiX6mvrqaznboI+8xFFayDqn2oeAh+bmuFaRtEUKS9XR9dvHTT6BrqotO6vB67ucaj0Ru6tn9zsB+xc6hqn2AInl+VWVEaJW8/VFgeZ6peoVWbCA6q90IW99L3AgejnYqJlR+ah5mFmoKZgpt7nXScdKJqp2Dq+ykY9woG+xD3V3KxcatwpBl+l3iXcpfPlL6irK0IrK6btr4asoGvd6wed6txomqYCJhqWpFLG/vR/WAG6vkRFfd2BsCygHWjH6R1l3BpGnSFdX53Hn54eXxzggiCcmqHXxv7XwYOc+DwFaRmrW63eAh4t8GCzBu+uZSesx+0nquloKwIoa2Wr7EasYGtd6ked6hto2Geb5hWmz6cPpxbnHmcCHicgqClGqiYpKWgHqCmtJbFG8K0f3SnH6h0m2mQXuaSGIm1gLF1rHWsbKRinAicY1yUVhtbX4N7ZB9jem1zd2wIdmuBamYaapNunHAenHGkdK15pn25fM18zHu2f56EqX+gfZh7CJh6knd1GnWEdn55Hn14d3xvgAiAb2uGZxtjZpKZax9qmnOdfKJ7ooGph68ygxiMW5hgpGUIDjv39hb5DPeA3/zLN/eA/QwHDqr4tvfDFTF8Tm5rHmxtWntFG2Npk5tvH2+bd6J/qAiAqYW4yhr4MSz8MgdAlE+dXx6dX6pqtXQIdLbCf84b0MKYprYftaWorpy1CJu1k8XSGvgyLAcOc/gPFves+WAFKgb7VfycfGR/ZIBkGYCvf7J8tftO+JwYJAb3qf1gBQ73kfe/Fvcr+LaRopKnlKwZjYCTb5he9yr8thjnBvdY+WAFLAb7BPxgfFB/V4JeGX7aeeBy5CT3/xj7Bgb7HPx4iH+AX3k/GYK8gLuAvPsA+GoYKQb3UP1gBQ5z9woW90r3jJKVlpyboxmUfJV9lXz3SfuTGPcIBvuf+Az3jPfoBSQG+yT7UnZueHF7chmAn3iocLH7F/dLGPsFBveI++z7qfwIBQ5z+AoW98MH97L4MQX7Awb7HvtnbFxwYXZmGXSzc7Nws/sh920Y+wYG96j8MQX7wwcOO/jeFt/8XQe2vvgm+IUF3/yUN/gjB3Rycm9xavwD/F8YNAcO+DoW5waAn4Sgh6EIiKCJv9wa9wkHsoqmiJoehaOCn36bfpt3mG+VCJZvZ5BfG15khX9pH2l+cXp5dHl1fm2DZuF/GJSwmqWfmQian6mStRu3rYF3oR+cfZNyZ4iLg38aaX9XgUODaYdxhnmHdIR2gnh+eH58en92CIB3hXNyGmCaZ6pwHm+qt33EG62skZapH6mXqp6sp45ykHaUeAhz93gVZIZugXgef3F4d3B8CHxxbYRpG2hxk5p6H3mbgp6jGpqPmZOXHpOYl5SakpqRpZGvkMuUu5armAgO9yfMFViuu3LIG8jAo7y3H7e7odDjGrGGroCsHoGrfad4o3mic51vmAiYbm2RaxtSW3RcZh/3lDP9YN0HtPgsFaynrJyxG7Gse2umH6ZrmFlHGkl9WW9qHmpvanplG1tmorhvH3qmg7jJGsqZvKesHg77U/f96BV2dG6AaRtgaJuqcB9wq3690RrQmb2nqh6rpq+buBuopIJ6oB+feZpxk2jgmBiBv3S0Z6cIqGddmVMbX2GBdmUfZnZua3lhCHhhglpUGjShSbZcHl22xHTSG8O7nKyyH7GtpLmUxjWXGIVffGt0dggO+HcW+WAz+5YHfKF3nHKYCJhzb5JsG2BlgHRoH2l1cWt6YQh6YYJcVxpWlVyeYh6eY6VrrnQIdK6xgLQby7ulvqwfSQf7g/gtFaumq5uzG7OsemqnH6ZqmVdEGkt+W3BsHmxwantkG2Vqm6xvH2+sfb3NGs+YvaWrHg74AuIVenRwgmsbX2eaqW4fbqp7tojECPgXBpWLk5Aa4XXNX7oeul9To0YbQ1FzW14fXlt1RzQaN6FKuFweXLfHdNcbx7yaqLIfsaimtJnAMJcYfmZ5cHR6CPtQ994VpqatmbMbuK96aacfnXWWa49fCPu1Bo64mq+npggO/DH3Qxb4V+/PJrsHqpCgl5YelpadkaYbm52JiJ0fmNgFkW1wjnIbZW2EfXYfdX19eIJ1CIV6iHFoGlQ9R9n8VwcO9Ps8FW+xvX3JG7+3lZ6uH6+fpaWbrQicrZPE3Br4VDpLB71jWaRNG15jgHRpH2l0cWt5YQh5YYJeWRpDnk6yVx5Ys8Jx0hvEu6K4sh9SiWWGeh6EbXx1dHoIe3Vsg2IbZW2Tm3YfepeBn4ilNpcYilOdYbFwCMX41RWrpqybsxuyrXtrqB+na5lbSxpJfVtwbB5sb2l7YxtiaZuqcB9wqn69zhrKmbqmqh4O9y4W968HtJCrlaIelKKcnaGZCJiio5KlG66mgXeeH553lGtfGvvc4/fcB76Fsn+mHn+ldqBvmgiab2qTZRtMWHNbYh/3ljP9YAcO/Gn3Lvj8Fe8zJwfj/PwV+Jsz/JsHDvtT9y4W92IHyMb3QfudBfcABvtu99r3WvdVBfsGBvtk+2cF+Cwz/WAHDvxp9ywW+WAz/WAHDvci9y4W96EHupCvlKQelaSanqCYCJigopKjG6yigXiZH5p3km5kGvvl4/fBB8GXsaOkHqOjqpevG6CchoKaH5qBln+QfAiRe45yaBr72+P3+AfGfbdvpx6ob2SZVxtJVW1OYh+BqHqhcpsIm3Nrk2UbaG2DfHAfcHt1d3tyCNQ8/JsHDvcuFvevB86ZuKaiHqOmq5ewG6OfhoCcH52Bl3ySegiSeY5wZxr7z+P30weziaiImx6GpIKhfp1+nXeacZYIlnFukWwbQ1RvUmUf1Tz8mwcO78YVXLjGdNMbubSWoLIfsaCoqJ+yCJ+xlb/OGt10y166HrpeUaJDG0tVeGReH1ZdcEQsGjOhSLhdHs738RWsqK+btxu3r3tqqB+oappaSxpHfFluah5qbmd6XxtfZ5usbh9urHy9zRrNmr2orB4O9y77WxX3kQeaeJ58on4If6Olhagbs7GWorAfr6GmrJ61CJ62lbrAGr2CuHq1Hnq0catqogiiaWSWXhtqboR+cx9zfnZ3eHEIzzv9Ygf3D/j0Fa6orJywG7Gre2qmH6ZqmVpJGkV9WG9qHmpwaXtkG2Vqm6twH3CrfrzNGs6ZvqiuHg74ePtbFfliPEUHwWdYpksbYmWAdmkfaXZxbHlhCHligVxXGjaiSLdaHlq3wHLJG6elkZijH6SYnpuYngj7kwf7e/j3Faymq5uxG7KsemioH6domVdGGkp+W3BsHmtwa3tlG2RqnKxvH26sfb3OGtCZvaWrHg77+vctFvejB7CQrZWrHpGflpualwiWmp2RnhugoIV/oR+q3AWebG2Ubht2eIV/eh96gHhyd2cI2jz8mwcO+1PuqhVvrr59zxu0r5KZqx+smaOfnKUInKWUpqkaqYSkfZ8efZ93mnOWcpVgmU2cYJZxk4KOfJGAk4SUCISVh5WWGp2Um5yYHpicqJKzG62lg3yeH558lnaPcOGXGIWtgaZ9n3yfdJttlgiXbGeRYxtwcYiEdB9zhHmCfYF5fnx7gXcIgHeGdnQacpFzmHYemHeeeqR/pH+3fcx7un+pgZiDCJyAlHt3GnWBeHh7Hnp3bYNjG2JslJ51H3WdfaaGrjR9GJVUoWKvbwgO/DH3b9YVfoGNj4QfhJCGkIiTCIiSiZukGvfE488z90kHM1YF+xRKR8z7vwdWj2mSeh6Se5d9nYEIgZykhqsbnqGOkKQff9gFiXt+ioIbDvh4FvibM/upB16GaoJzHoF0e3l0fQh+dHKEcRtwdZKYeR96mH+dhaIIiJuJqrka97Mz+9UHZY1wjnoekXGUdZd6mHmffKWACH+mp4WqG9DCqMazHz4HDvtT97gW91n4mwUxBvsI+9F9ZYBqhHAZgK+Arn+s+wP3yxgtBvdY/JsFDqr3kRb0+COfM977ywXmBvc3+JsFNQYx+8BuJ3HuPffBBTEGOfvEekmCaIqFGW33BDj3vwUwBvcw/JsFDvtT9wUW9x/3WqRl9vs0BfYG+1D3ofdE944FIAY1+w5/en54fHYZgpp/nnyhOfcPGPsABvdE+477UvuhBQ77U/cL+2YVp6OSmJ8foJmdoJqol6CbsqHE91j4pBgzBvsD+8N9ZX9kgWQZgLR+s32x+wD3wBgtBvdZ/J2HgomEiYYZf2iCdYWChH+Bgn+FCISAe4h3G316jpB4H5U6BYSgnoecGw77U/hzFtf7hQdpZomIYx/ByPeu990Fxfw7RPdmB6esjI2wH/vc/A8FQwcO+L33dBXS/L9EBw6Liwb4wBT5RxUAAAMCJAH0AAUAAAKKArsAAACMAooCuwAAAd8AMQECAAAAAAYAAAAAAAAAgAAAARAAAAAAAAAAAAAAACoyMSoAAAAg4AAD7v67AGQD7gFFAAAAAAAAAAACBwLMAAAAIAADAAAAAQADAAEAAAAMAAQAcAAAABgAEAADAAgAIAApACsALgA5AEkAWgBpAHogE+AA//8AAAAgACgAKwAuADAAQQBLAGEAayAT4AD////h/9r/2f/X/9b/z//O/8j/x+AvIAEAAQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABAAAAABAAAAAAAF8PPPUAAAPoAAAAAJ4LficAAAAAngt+JwAA/rsP/wPuAAAAEQAAAAAAAAAAAAEAAAPu/rsAAP//AAAAAAAAAswAAAAAAAAAAAAAAAAAAABDAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAB8AAAAfAAAAAAAAAAAAAABXAAAAHwAAAAAAAAAAAAAAAAAAAI4AAAAfAAAAVwAAAAAAAABXAAAAHwAAAAAAAAAAAAAAHwAAAAAAAAD9AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAACOAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAHwAAAAAAAAAAAAAAAAAAAAAAAAAAUAAAQwAAAAAAFAD2AAEAAAAAAAAAEAAAAAEAAAAAAAEADgAQAAEAAAAAAAIABwAeAAEAAAAAAAMACAAlAAEAAAAAAAQADgAtAAEAAAAAAAUADAA7AAEAAAAAAAYAAABHAAEAAAAAAAcABwBHAAEAAAAAAAgABwBOAAEAAAAAAAkABwBVAAMAAQQJAAAAIABcAAMAAQQJAAEAHAB8AAMAAQQJAAIADgCYAAMAAQQJAAMAEACmAAMAAQQJAAQAHAC2AAMAAQQJAAUAGADSAAMAAQQJAAYAAADqAAMAAQQJAAcADgDqAAMAAQQJAAgADgD4AAMAAQQJAAkADgEGT3JpZ2luYWwgbGljZW5jZUJPR0JERCtBcmlhbE1UVW5rbm93bnVuaXF1ZUlEQk9HQkREK0FyaWFsTVRWZXJzaW9uIDAuMTFVbmtub3duVW5rbm93blVua25vd24ATwByAGkAZwBpAG4AYQBsACAAbABpAGMAZQBuAGMAZQBCAE8ARwBCAEQARAArAEEAcgBpAGEAbABNAFQAVQBuAGsAbgBvAHcAbgB1AG4AaQBxAHUAZQBJAEQAQgBPAEcAQgBEAEQAKwBBAHIAaQBhAGwATQBUAFYAZQByAHMAaQBvAG4AIAAwAC4AMQAxAFUAbgBrAG4AbwB3AG4AVQBuAGsAbgBvAHcAbgBVAG4AawBuAG8AdwBuAAAAAwAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA==); }&#xA;@font-face { font-family: &quot;g_font_9&quot;; src: url(data:font/opentype;base64,AAEAAAANAIAAAwBQT1MvMrStPVsAAADcAAAAYGNtYXBG2wq5AAABPAAAGuxjdnQgoRzX6wAAHCgAAAZUZnBnbcx5WZoAACJ8AAAGbmdseWYGJQCaAAAo7AAAAGJoZWFk53kpCAAAKVAAAAA2aGhlYRIzFiYAACmIAAAAJGhtdHh0wP1UAAAprAAANXRsb2NhAATFOgAAXyAAADV4bWF4cBK5AcEAAJSYAAAAIG5hbWXjLEesAACUuAAAAf5wb3N0AAMAAAAAlrgAAAAgcHJlcCXWTb8AAJbYAAALvgADAiQB9AAFAAACigK7AAAAjAKKArsAAAHfADEBAgAAAAAGAAAAAAAAAAAAAAAQACAAAAAAAAAAAAAqMjEqAAAlz+1bBz7+TgBkCAwCmQAAAAAAAAAAAgMCzgAAJc8AAwAAAAEAAwABAAAADAAEGuAAAAAGAAQAAQACJc/tW///AAAlz+AA///bxQAAAAEAAAAEAAAAAAABAAIAAwAEAAUABgAHAAgACQAKAAsADAANAA4ADwAQABEAEgATABQAFQAWABcAGAAZABoAGwAcAB0AHgAfACAAIQAiACMAJAAlACYAJwAoACkAKgArACwALQAuAC8AMAAxADIAMwA0ADUANgA3ADgAOQA6ADsAPAA9AD4APwBAAEEAQgBDAEQARQBGAEcASABJAEoASwBMAE0ATgBPAFAAUQBSAFMAVABVAFYAVwBYAFkAWgBbAFwAXQBeAF8AYABhAGIAYwBkAGUAZgBnAGgAaQBqAGsAbABtAG4AbwBwAHEAcgBzAHQAdQB2AHcAeAB5AHoAewB8AH0AfgB/AIAAgQCCAIMAhACFAIYAhwCIAIkAigCLAIwAjQCOAI8AkACRAJIAkwCUAJUAlgCXAJgAmQCaAJsAnACdAJ4AnwCgAKEAogCjAKQApQCmAKcAqACpAKoAqwCsAK0ArgCvALAAsQCyALMAtAC1ALYAtwC4ALkAugC7ALwAvQC+AL8AwADBAMIAwwDEAMUAxgDHAMgAyQDKAMsAzADNAM4AzwDQANEA0gDTANQA1QDWANcA2ADZANoA2wDcAN0A3gDfAOAA4QDiAOMA5ADlAOYA5wDoAOkA6gDrAOwA7QDuAO8A8ADxAPIA8wD0APUA9gD3APgA+QD6APsA/AD9AP4A/wEAAQEBAgEDAQQBBQEGAQcBCAEJAQoBCwEMAQ0BDgEPARABEQESARMBFAEVARYBFwEYARkBGgEbARwBHQEeAR8BIAEhASIBIwEkASUBJgEnASgBKQEqASsBLAEtAS4BLwEwATEBMgEzATQBNQE2ATcBOAE5AToBOwE8AT0BPgE/AUABQQFCAUMBRAFFAUYBRwFIAUkBSgFLAUwBTQFOAU8BUAFRAVIBUwFUAVUBVgFXAVgBWQFaAVsBXAFdAV4BXwFgAWEBYgFjAWQBZQFmAWcBaAFpAWoBawFsAW0BbgFvAXABcQFyAXMBdAF1AXYBdwF4AXkBegF7AXwBfQF+AX8BgAGBAYIBgwGEAYUBhgGHAYgBiQGKAYsBjAGNAY4BjwGQAZEBkgGTAZUBlgGXAZgBmQGaAZsBnAGdAZ4BnwGgAaEBogGjAaQBpQGmAacBqAGpAaoBqwGsAa0BrgGvAbABsQGyAbMBtAG1AbYBtwG4AbkBugG7AbwBvQG+Ab8BwAHBAcIBwwHEAcUBxgHHAcgByQHKAcsBzAHNAc4BzwHQAdEB0gHTAdQB1QHWAdcB2AHZAdoB2wHcAd0B3gHfAeAB4QHiAeMB5AHlAeYB5wHoAekB6gHrAewB7QHuAe8B8AHxAfIB8wH0AfUB9gH3AfgB+QH6AfsB/AH9Af4B/wIAAgECAgIDAgQCBQIGAgcCCAIJAgoCCwIMAg0CDgIPAhACEQISAhMCFAIVAhYCFwIYAhkCGgIbAhwCHQIeAh8CIAIhAiICIwIkAiUCJgInAigCKQIqAisCLAItAi4CLwIwAjECMgIzAjQCNQI2AjcCOAI5AjoCOwI8Aj0CPgI/AkACQQJCAkMCRAJFAkYCRwJIAkkCSgJLAkwCTQJOAk8CUAJRAlICUwJUAlUCVgJXAlgCWQJaAlsCXAJdAl4CXwJgAmECYgJjAmQCZQJmAmcCaAJpAmoCawJsAm0CbgJvAnACcQJyAnMCdAJ1AnYCdwJ4AnkCegJ7AnwCfQJ+An8CgAKBAoICgwKEAoUChgKHAogCiQKKAosCjAKNAo4CjwKQApECkgKTApQClQKWApcCmAKZApoCmwKcAp0CngKfAqACoQKiAqMCpAKlAqYCpwKoAqkCqgKrAqwCrQKuAq8CsAKxArICswK0ArUCtgK3ArgCuQK6ArsCvAK9Ar4CvwLAAsECwgLDAsQCxQLGAscCyALJAsoCywLMAs0CzgLPAtAC0QLSAtMC1ALVAtYC1wLYAtkC2gLbAtwC3QLeAt8C4ALhAuIC4wLkAuUC5gLnAugC6QLqAusC7ALtAu4C7wLwAvEC8gLzAvQC9QL2AvcC+AL5AvoC+wL8Av0C/gL/AwADAQMCAwMDBAMFAwYDBwMIAwkDCgMLAwwDDQMOAw8DEAMRAxIDEwMUAxUDFgMXAxgDGQMaAxsDHAMdAx4DHwMgAyEDIgMjAyQDJQMmAycDKAMpAyoDKwMsAy0DLgMvAzADMQMyAzMDNAM1AzYDNwM4AzkDOgM7AzwDPQM+Az8DQANBA0IDQwNEA0UDRgNHA0gDSQNKA0sDTANNA04DTwNQA1EDUgNTA1QDVQNWA1cDWANZA1oDWwNcA10DXgNfA2ADYQNiA2MDZANlA2YDZwNoA2kDagNrA2wDbQNuA28DcANxA3IDcwN0A3UDdgN3A3gDeQN6A3sDfAN9A34DfwOAA4EDggODA4QDhQOGA4cDiAOJA4oDiwOMA40DjgOPA5ADkQOSA5MDlAOVA5YDlwOYA5kDmgObA5wDnQOeA58DoAOhA6IDowOkA6UDpgOnA6gDqQOqA6sDrAOtA64DrwOwA7EDsgOzA7QDtQO2A7cDuAO5A7oDuwO8A70DvgO/A8ADwQPCA8MDxAPFA8YDxwPIA8kDygPLA8wDzQPOA88D0APRA9ID0wPUA9UD1gPXA9gD2QPaA9sD3APdA94D3wPgA+ED4gPjA+QD5QPmA+cD6APpA+oD6wPsA+0D7gPvA/AD8QPyA/MD9AP1A/YD9wP4A/kD+gP7A/wD/QP+A/8EAAQBBAIEAwQEBAUEBgQHBAgECQQKBAsEDAQNBA4EDwQQBBEEEgQTBBQEFQQWBBcEGAQZBBoEGwQcBB0EHgQfBCAEIQQiBCMEJAQlBCYEJwQoBCkEKgQrBCwELQQuBC8EMAQxBDIEMwQ0BDUENgQ3BDgEOQQ6BDsEPAQ9BD4EPwRABEEEQgRDBEQERQRGBEcESARJBEoESwRMBE0ETgRPBFAEUQRSBFMEVARVBFYEVwRYBFkEWgRbBFwEXQReBF8EYARhBGIEYwRkBGUEZgRnBGgEaQRqBGsEbARtBG4EbwRwBHEEcgRzBHQEdQR2BHcEeAR5BHoEewR8BH0EfgR/BIAEgQSCBIMEhASFBIYEhwSIBIkEigSLBIwEjQSOBI8EkASRBJIEkwSUBJUElgSXBJgEmQSaBJsEnASdBJ4EnwSgBKEEogSjBKQEpQSmBKcEqASpBKoEqwSsBK0ErgSvBLAEsQSyBLMEtAS1BLYEtwS4BLkEugS7BLwEvQS+BL8EwATBBMIEwwTEBMUExgTHBMgEyQTKBMsEzATNBM4EzwTQBNEE0gTTBNQE1QTWBNcE2ATZBNoE2wTcBN0E3gTfBOAE4QTiBOME5ATlBOYE5wToBOkE6gTrBOwE7QTuBO8E8ATxBPIE8wT0BPUE9gT3BPgE+QT6BPsE/AT9BP4E/wUABQEFAgUDBQQFBQUGBQcFCAUJBQoFCwUMBQ0FDgUPBRAFEQUSBRMFFAUVBRYFFwUYBRkFGgUbBRwFHQUeBR8FIAUhBSIFIwUkBSUFJgUnBSgFKQUqBSsFLAUtBS4FLwUwBTEFMgUzBTQFNQU2BTcFOAU5BToFOwU8BT0FPgU/BUAFQQVCBUMFRAVFBUYFRwVIBUkFSgVLBUwFTQVOBU8FUAVRBVIFUwVUBVUFVgVXBVgFWQVaBVsFXAVdBV4FXwVgBWEFYgVjBWQFZQVmBWcFaAVpBWoFawVsBW0FbgVvBXAFcQVyBXMFdAV1BXYFdwV4BXkFegV7BXwFfQV+BX8FgAWBBYIFgwWEBYUFhgWHBYgFiQWKBYsFjAWNBY4FjwWQBZEFkgWTBZQFlQWWBZcFmAWZBZoFmwWcBZ0FngWfBaAFoQWiBaMFpAWlBaYFpwWoBakFqgWrBawFrQWuBa8FsAWxBbIFswW0BbUFtgW3BbgFuQW6BbsFvAW9Bb4FvwXABcEFwgXDBcQFxQXGBccFyAXJBcoFywXMBc0FzgXPBdAF0QXSBdMF1AXVBdYF1wXYBdkF2gXbBdwF3QXeBd8F4AXhBeIF4wXkBeUF5gXnBegF6QXqBesF7AXtBe4F7wXwBfEF8gXzBfQF9QX2BfcF+AX5BfoF+wX8Bf0F/gX/BgAGAQYCBgMGBAYFBgYGBwYIBgkGCgYLBgwGDQYOBg8GEAYRBhIGEwYUBhUGFgYXBhgGGQYaBhsGHAYdBh4GHwYgBiEGIgYjBiQGJQYmBicGKAYpBioGKwYsBi0GLgYvBjAGMQYyBjMGNAY1BjYGNwY4BjkGOgY7BjwGPQY+Bj8GQAZBBkIGQwZEBkUGRgZHBkgGSQZKBksGTAZNBk4GTwZQBlEGUgZTBlQGVQZWBlcGWAZZBloGWwZcBl0GXgZfBmAGYQZiBmMGZAZlBmYGZwZoBmkGagZrBmwGbQZuBm8GcAZxBnIGcwZ0BnUGdgZ3BngGeQZ6BnsGfAZ9Bn4GfwaABoEGggaDBoQGhQaGBocGiAaJBooGiwaMBo0GjgaPBpAGkQaSBpMGlAaVBpYGlwaYBpkGmgabBpwGnQaeBp8GoAahBqIGowakBqUGpganBqgGqQaqBqsGrAatBq4GrwawBrEGsgazBrQGtQa2BrcGuAa5BroGuwa8Br0Gvga/BsAGwQbCBsMGxAbFBsYGxwbIBskGygbLBswGzQbOBs8G0AbRBtIG0wbUBtUG1gbXBtgG2QbaBtsG3AbdBt4G3wbgBuEG4gbjBuQG5QbmBucG6AbpBuoG6wbsBu0G7gbvBvAG8QbyBvMG9Ab1BvYG9wb4BvkG+gb7BvwG/Qb+Bv8HAAcBBwIHAwcEBwUHBgcHBwgHCQcKBwsHDAcNBw4HDwcQBxEHEgcTBxQHFQcWBxcHGAcZBxoHGwccBx0HHgcfByAHIQciByMHJAclByYHJwcoBykHKgcrBywHLQcuBy8HMAcxBzIHMwc0BzUHNgc3BzgHOQc6BzsHPAc9Bz4HPwdAB0EHQgdDB0QHRQdGB0cHSAdJB0oHSwdMB00HTgdPB1AHUQdSB1MHVAdVB1YHVwdYB1kHWgdbB1wHXQdeB18HYAdhB2IHYwdkB2UHZgdnB2gHaQdqB2sHbAdtB24HbwdwB3EHcgdzB3QHdQd2B3cHeAd5B3oHewd8B30Hfgd/B4AHgQeCB4MHhAeFB4YHhweIB4kHigeLB4wHjQeOB48HkAeRB5IHkweUB5UHlgeXB5gHmQeaB5sHnAedB54HnwegB6EHogejB6QHpQemB6cHqAepB6oHqwesB60HrgevB7AHsQeyB7MHtAe1B7YHtwe4B7kHuge7B7wHvQe+B78HwAfBB8IHwwfEB8UHxgfHB8gHyQfKB8sHzAfNB84HzwfQB9EH0gfTB9QH1QfWB9cH2AfZB9oH2wfcB90H3gffB+AH4QfiB+MH5AflB+YH5wfoB+kH6gfrB+wH7QfuB+8H8AfxB/IH8wf0B/UH9gf3B/gH+Qf6B/sH/Af9B/4H/wgACAEIAggDCAQIBQgGCAcICAgJCAoICwgMCA0IDggPCBAIEQgSCBMIFAgVCBYIFwgYCBkIGggbCBwIHQgeCB8IIAghCCIIIwgkCCUIJggnCCgIKQgqCCsILAgtCC4ILwgwCDEIMggzCDQINQg2CDcIOAg5CDoIOwg8CD0IPgg/CEAIQQhCCEMIRAhFCEYIRwhICEkISghLCEwITQhOCE8IUAhRCFIIUwhUCFUIVghXCFgIWQhaCFsIXAhdCF4IXwhgCGEIYghjCGQIZQhmCGcIaAhpCGoIawhsCG0IbghvCHAIcQhyCHMIdAh1CHYIdwh4CHkIegh7CHwIfQh+CH8IgAiBCIIIgwiECIUIhgiHCIgIiQiKCIsIjAiNCI4IjwiQCJEIkgiTCJQIlQiWCJcImAiZCJoImwicCJ0IngifCKAIoQiiCKMIpAilCKYIpwioCKkIqgirCKwIrQiuCK8IsAixCLIIswi0CLUItgi3CLgIuQi6CLsIvAi9CL4IvwjACMEIwgjDCMQIxQjGCMcIyAjJCMoIywjMCM0IzgjPCNAI0QjSCNMI1AjVCNYI1wjYCNkI2gjbCNwI3QjeCN8I4AjhCOII4wjkCOUI5gjnCOgI6QjqCOsI7AjtCO4I7wjwCPEI8gjzCPQI9Qj2CPcI+Aj5CPoI+wj8CP0I/gj/CQAJAQkCCQMJBAkFCQYJBwkICQkJCgkLCQwJDQkOCQ8JEAkRCRIJEwkUCRUJFgkXCRgJGQkaCRsJHAkdCR4JHwkgCSEJIgkjCSQJJQkmCScJKAkpCSoJKwksCS0JLgkvCTAJMQkyCTMJNAk1CTYJNwk4CTkJOgk7CTwJPQk+CT8JQAlBCUIJQwlECUUJRglHCUgJSQlKCUsJTAlNCU4JTwlQCVEJUglTCVQJVQlWCVcJWAlZCVoJWwlcCV0JXglfCWAJYQliCWMJZAllCWYJZwloCWkJaglrCWwJbQluCW8JcAlxCXIJcwl0CXUJdgl3CXgJeQl6CXsJfAl9CX4JfwmACYEJggmDCYQJhQmGCYcJiAmJCYoJiwmMCY0JjgmPCZAJkQmSCZMJlAmVCZYJlwmYCZkJmgmbCZwJnQmeCZ8JoAmhCaIJowmkCaUJpgmnCagJqQmqCasJrAmtCa4JrwmwCbEJsgmzCbQJtQm2CbcJuAm5CboJuwm8Cb0Jvgm/CcAJwQnCCcMJxAnFCcYJxwnICckJygnLCcwJzQnOCc8J0AnRCdIJ0wnUCdUJ1gnXCdgJ2QnaCdsJ3AndCd4J3wngCeEJ4gnjCeQJ5QnmCecJ6AnpCeoJ6wnsCe0J7gnvCfAJ8QnyCfMJ9An1CfYJ9wn4CfkJ+gn7CfwJ/Qn+Cf8KAAoBCgIKAwoECgUKBgoHCggKCQoKCgsKDAoNCg4KDwoQChEKEgoTChQKFQoWChcKGAoZChoKGwocCh0KHgofCiAKIQoiCiMKJAolCiYKJwooCikKKgorCiwKLQouCi8KMAoxCjIKMwo0CjUKNgo3CjgKOQo6CjsKPAo9Cj4KPwpACkEKQgpDCkQKRQpGCkcKSApJCkoKSwpMCk0KTgpPClAKUQpSClMKVApVClYKVwpYClkKWgpbClwKXQpeCl8KYAphCmIKYwpkCmUKZgpnCmgKaQpqCmsKbAptCm4KbwpwCnEKcgpzCnQKdQp2CncKeAp5CnoKewp8Cn0Kfgp/CoAKgQqCCoMKhAqFCoYKhwqICokKigqLCowKjQqOCo8KkAqRCpIKkwqUCpUKlgqXCpgKmQqaCpsKnAqdCp4KnwqgCqEKogqjCqQKpQqmCqcKqAqpCqoKqwqsCq0KrgqvCrAKsQqyCrMKtAq1CrYKtwq4CrkKugq7CrwKvQq+Cr8KwArBCsIKwwrECsUKxgrHCsgKyQrKCssKzArNCs4KzwrQCtEK0grTCtQK1QrWCtcK2ArZCtoK2wrcCt0K3grfCuAK4QriCuMK5ArlCuYK5wroCukK6grrCuwK7QruCu8K8ArxCvIK8wr0CvUK9gr3CvgK+Qr6CvsK/Ar9Cv4K/wsACwELAgsDCwQLBQsGCwcLCAsJCwoLCwsMCw0LDgsPCxALEQsSCxMLFAsVCxYLFwsYCxkLGgsbCxwLHQseCx8LIAshCyILIwskCyULJgsnCygLKQsqCysLLAstCy4LLwswCzELMgszCzQLNQs2CzcLOAs5CzoLOws8Cz0LPgs/C0ALQQtCC0MLRAtFC0YLRwtIC0kLSgtLC0wLTQtOC08LUAtRC1ILUwtUC1ULVgtXC1gLWQtaC1sLXAtdC14LXwtgC2ELYgtjC2QLZQtmC2cLaAtpC2oLawtsC20LbgtvC3ALcQtyC3MLdAt1C3YLdwt4C3kLegt7C3wLfQt+C38LgAuBC4ILgwuEC4ULhguHC4gLiQuKC4sLjAuNC44LjwuQC5ELkguTC5QLlQuWC5cLmAuZC5oLmwucC50LngufC6ALoQuiC6MLpAulC6YLpwuoC6kLqgurC6wLrQuuC68LsAuxC7ILswu0C7ULtgu3C7gLuQu6C7sLvAu9C74LvwvAC8ELwgvDC8QLxQvGC8cLyAvJC8oLywvMC80LzgvPC9AL0QvSC9ML1AvVC9YL1wvYC9kL2gvbC9wL3QveC98L4AvhC+IL4wvkC+UL5gvnC+gL6QvqC+sL7AvtC+4L7wvwC/EL8gvzC/QL9Qv2C/cL+Av5C/oL+wv8C/0L/gv/DAAMAQwCDAMMBAwFDAYMBwwIDAkMCgwLDAwMDQwODA8MEAwRDBIMEwwUDBUMFgwXDBgMGQwaDBsMHAwdDB4MHwwgDCEMIgwjDCQMJQwmDCcMKAwpDCoMKwwsDC0MLgwvDDAMMQwyDDMMNAw1DDYMNww4DDkMOgw7DDwMPQw+DD8MQAxBDEIMQwxEDEUMRgxHDEgMSQxKDEsMTAxNDE4MTwxQDFEMUgxTDFQMVQxWDFcMWAxZDFoMWwxcDF0MXgxfDGAMYQxiDGMMZAxlDGYMZwxoDGkMagxrDGwMbQxuDG8McAxxDHIMcwx0DHUMdgx3DHgMeQx6DHsMfAx9DH4MfwyADIEMggyDDIQMhQyGDIcMiAyJDIoMiwyMDI0MjgyPDJAMkQySDJMMlAyVDJYMlwyYDJkMmgybDJwMnQyeDJ8MoAyhDKIMowykDKUMpgynDKgMqQyqDKsMrAytDK4MrwywDLEMsgyzDLQMtQy2DLcMuAy5DLoMuwy8DL0Mvgy/DMAMwQzCDMMMxAzFDMYMxwzIDMkMygzLDMwMzQzODM8M0AzRDNIM0wzUDNUM1gzXDNgM2QzaDNsM3AzdDN4M3wzgDOEM4gzjDOQM5QzmDOcM6AzpDOoM6wzsDO0M7gzvDPAM8QzyDPMM9Az1DPYM9wz4DPkM+gz7DPwM/Qz+DP8NAA0BDQINAw0EDQUNBg0HDQgNCQ0KDQsNDA0NDQ4NDw0QDRENEg0TDRQNFQ0WDRcNGA0ZDRoNGw0cDR0NHg0fDSANIQ0iDSMNJA0lDSYNJw0oDSkNKg0rDSwNLQ0uDS8NMA0xDTINMw00DTUNNg03DTgNOQ06DTsNPA09DT4NPw1ADUENQg1DDUQNRQ1GDUcNSA1JDUoNSw1MDU0NTg1PDVANUQ1SDVMNVA1VDVYNVw1YDVkNWg1bDVwFugAZBboAGgWnABkEJgAYAAD/5wAA/+gAAP/n/mn/6AW6ABn+af/oAuoAAAC4AAAAuAAAAAAAqACtAWkArQC/AMIB8AAYAK8AuQC0AMgAFwBEAJwAfACUAIcABgBaAMgAiQBSAFIABQBEAJQBGf+0AC8AoQADAKEAzQAXAFcAfgC6ABYBGP/pAH8AhQPTAIcAhQANACIAQQBQAG8AjQFM/3UAXADfBIMANwBMAG4AcAGA/1j/jv+S/6QApQC5A8j//QALABoAYwBjAM3/7gXY/9wALQBcAJUAmQDfAZIJtQBAAFcAgAC5A50AcgCaA10EAf9n//oAAwAhAHcAzQAEAE0AzQHAAisATABlAOcBGAF8A0MF2P+j/7D/xAADABwAXQBoAJoAugE1AUcCIQVc/03/zQAWAC0AeACAAJkAsgC2ALYAuAC9ANoBDAXw/6T/8AAZACwASQB/ALQAzgHAA/79gf4/AAAABQAYACkAOQBJAG8AvgDHANABIwHBAm8FDAUyBUAFev/UABQAMQBVAFcApwC0AOYB9wJ+An4CfwPGBEb/QgAOAIUAkQC/AMIAxQDhARoBLwFPAVYCKQJvAp4DcgAIACwAMQAxAGQAaQCJAJgAxwDeASsBtgIMAs8DowSrBPsGHf7g/w4ABgAmAJsAnQDBAQ0BGAEgAXMBggHWAeMCQwJfApsC4gOUBKkE0gdhABwAXgBtAI0AqwD3ARIBOAFRAVsBaAF8AYcBkQGZAc0B0AHoAkECVAJrAu8DaANxA70EQgRCBFMEcwSDBYYFiwbo/lj+xP7R/vf/Mv+GAFEAfACBAJEAlQCeALQAuQDPANkA2QDfAOIBBQELAQ4BDgEgASEBVQF7AXsBfgGNAaIBqAGpAbQB0AHQAeIB6QHyAfUB+wIAAgACBgIbAiECIgIiAiMCcgJ3ApQCnALPAs8C0ALsAvkDFwMiAysDNQM8A1kDbwNxA4cDkAOQA7UD4QQaBM8E/wUyBTIFlgWfBagFqwXCBfAGDAeCCAAIzPyj/Sr93v4A/oj+lv6y/rT/4QAVABkAGgAcAB8APABRAGEAYQBqAHgAlgClAK8A0wEMARgBGgEqAT4BTAFRAV8BagFxAXgBggGEAZoBpQGoAakBrgG8Ac0B1wHvAgACDQIcAiECIgIuAjUCQgJPAk8CXgJlAnECkAKSArQC1gL6AwcDCwMPAxUDKgNHA10DZQN0A3kDlgOwA8wD3QPiA/YD/AP8A/8ECgQfBCIEJgQrBEcEXwR1BJ4E5wTnBVwFywXlBgoGbQaGBrgG8Qc2Bz4HUAdRB10Hjwe2B9QIYAC2AMMAtQC3AAAAAAAAAAAAAAAAAeADgQNFA7UAjgIzBBkCzgLOAC0AXwBkA00CPwAAAqgBiAJ9AbQCJAV4BjsCOwFOAPAEJgKUAsYCnwL2AjsDTQFLAVMAagIxAAAAAAAABhQEqgAAADwEwwDtBLwCZQLOA7UAeAYMAX4C7wYMALIBAAI5AAABxQMwBCsDywDaA98BBwShANsECgEXAe0CpwNQAQsBvQQ+BVgAIQOcAK4DcQF9ALUCRQAACvsIjAErAU4BqgCHAFQBMgH4A/8AAwJOALQANwPjAIMAawLYAO0AdwCIAJcBZARnAI4AMwF8AOcApgKeAykFbgYqBhUByQJpBIoCEwG0AAIEqQAAAjkBJAEDBRQAhAFdA5oG7wLZAHUAzwQKAN4DrAS8As8CrgNNBPAFUgFoAG0AfQCGAHH/gQB5BVgE0gFnAAMBVgAlBOAAlAB8AzIEIQCUAH8AcgBcAC8AtgAYALoAuABBA00AcgAYAB8ATAFqAVUAmQCaAJoAmACyAAQAeABpABQAVwBuAM4AtAZUArgAZwUOAWUA5wAABMv+UgBa/6YAmf9nAG7/kgAt/9QAh/98ALgAqADlAI8AqAGF/nsAcAAeANkA3gFMBUYCzwVG/y0CigLZAlMClgC3AAAAAAAAAAAAAAAAAAABJQEYAOoA6gCuAAAAPgW7AIoE1wBTAD//jP/VABUAKAAiAJkAYgBKAOQAbQDuAOUASAPAADP+TgKx/0YDcAB5Bd8AUf+n/x8BCgBo/2wATwC8AKUHBQBhBysA7QSwAdIAtgB7AGUCUv90A2X+aQCUAI8AXABAAIYAdQCJAIlAQ1VUQUA/Pj08Ozo5ODc1NDMyMTAvLi0sKyopKCcmJSQjIiEgHx4dHBsaGRgXFhUUExIREA8ODQwLCgkIBwYFBAMCAQAsRSNGYCCwJmCwBCYjSEgtLEUjRiNhILAmYbAEJiNISC0sRSNGYLAgYSCwRmCwBCYjSEgtLEUjRiNhsCBgILAmYbAgYbAEJiNISC0sRSNGYLBAYSCwZmCwBCYjSEgtLEUjRiNhsEBgILAmYbBAYbAEJiNISC0sARAgPAA8LSwgRSMgsM1EIyC4AVpRWCMgsI1EI1kgsO1RWCMgsE1EI1kgsJBRWCMgsA1EI1khIS0sICBFGGhEILABYCBFsEZ2aIpFYEQtLAGxCwpDI0NlCi0sALEKC0MjQwstLACwFyNwsQEXPgGwFyNwsQIXRTqxAgAIDS0sRbAaI0RFsBkjRC0sIEWwAyVFYWSwUFFYRUQbISFZLSywAUNjI2KwACNCsA8rLSwgRbAAQ2BELSwBsAZDsAdDZQotLCBpsEBhsACLILEswIqMuBAAYmArDGQjZGFcWLADYVktLEWwESuwFyNEsBd65BgtLEWwESuwFyNELSywEkNYh0WwESuwFyNEsBd65BsDikUYaSCwFyNEioqHILCgUViwESuwFyNEsBd65BshsBd65FlZGC0sLSywAiVGYIpGsEBhjEgtLEtTIFxYsAKFWViwAYVZLSwgsAMlRbAZI0RFsBojREVlI0UgsAMlYGogsAkjQiNoimpgYSCwGoqwAFJ5IbIaGkC5/+AAGkUgilRYIyGwPxsjWWFEHLEUAIpSebMZQCAZRSCKVFgjIbA/GyNZYUQtLLEQEUMjQwstLLEOD0MjQwstLLEMDUMjQwstLLEMDUMjQ2ULLSyxDg9DI0NlCy0ssRARQyNDZQstLEtSWEVEGyEhWS0sASCwAyUjSbBAYLAgYyCwAFJYI7ACJTgjsAIlZTgAimM4GyEhISEhWQEtLEuwZFFYRWmwCUNgihA6GyEhIVktLAGwBSUQIyCK9QCwAWAj7ewtLAGwBSUQIyCK9QCwAWEj7ewtLAGwBiUQ9QDt7C0sILABYAEQIDwAPC0sILABYQEQIDwAPC0ssCsrsCoqLSwAsAdDsAZDCy0sPrAqKi0sNS0sdrgCIyNwECC4AiNFILAAUFiwAWFZOi8YLSwhIQxkI2SLuEAAYi0sIbCAUVgMZCNki7ggAGIbsgBALytZsAJgLSwhsMBRWAxkI2SLuBVVYhuyAIAvK1mwAmAtLAxkI2SLuEAAYmAjIS0stAABAAAAFbAIJrAIJrAIJrAIJg8QFhNFaDqwARYtLLQAAQAAABWwCCawCCawCCawCCYPEBYTRWhlOrABFi0sS1MjS1FaWCBFimBEGyEhWS0sS1RYIEWKYEQbISFZLSxLUyNLUVpYOBshIVktLEtUWDgbISFZLSywE0NYAxsCWS0ssBNDWAIbA1ktLEtUsBJDXFpYOBshIVktLLASQ1xYDLAEJbAEJQYMZCNkYWS4BwhRWLAEJbAEJQEgRrAQYEggRrAQYEhZCiEhGyEhWS0ssBJDXFgMsAQlsAQlBgxkI2RhZLgHCFFYsAQlsAQlASBGuP/wYEggRrj/8GBIWQohIRshIVktLEtTI0tRWliwOisbISFZLSxLUyNLUVpYsDsrGyEhWS0sS1MjS1FasBJDXFpYOBshIVktLAyKA0tUsAQmAktUWoqKCrASQ1xaWDgbISFZLSxLUliwBCWwBCVJsAQlsAQlSWEgsABUWCEgQ7AAVViwAyWwAyW4/8A4uP/AOFkbsEBUWCBDsABUWLACJbj/wDhZGyBDsABUWLADJbADJbj/wDi4/8A4G7ADJbj/wDhZWVlZISEhIS0sRiNGYIqKRiMgRopgimG4/4BiIyAQI4q5AsICwopwRWAgsABQWLABYbj/uosbsEaMWbAQYGgBOi0ssQIAQrEjAYhRsUABiFNaWLkQAAAgiFRYsgIBAkNgQlmxJAGIUVi5IAAAQIhUWLICAgJDYEKxJAGIVFiyAiACQ2BCAEsBS1JYsgIIAkNgQlkbuUAAAICIVFiyAgQCQ2BCWblAAACAY7gBAIhUWLICCAJDYEJZuUAAAQBjuAIAiFRYsgIQAkNgQlm5QAACAGO4BACIVFiyAkACQ2BCWVlZWVktLLACQ1RYS1MjS1FaWDgbISFZGyEhISFZLQAAAAIBAAAABQAFAAADAAcAACERIRElIREhAQAEAPwgA8D8QAUA+wAgBMAAAAEAsgCJBCMD+gANAAABMhYWFRQAIyIANTQ2NgJrbtR2/v62t/7+dtQD+nLUcrf+/gECt3PTcgAAAAABAAAABThSAAAAAF8PPPUIOwgAAAAAAKLjJyoAAAAA0pR/Gvqv/WcQAAgMAAAACQABAAEAAAAAAAEAAAc+/k4AQxAA+q/6ehAAAAEAAAAAAAAAAAAAAAAAAA1dBgABAAAAAAACOQAAAjkAAAI5ALAC1wBeBHMAFQRzAEkHHQB3BVYAWAGHAFoCqgB8AqoAfAMdAEAErAByAjkAqgKqAEECOQC6AjkAAARzAFUEcwDfBHMAPARzAFYEcwAaBHMAVQRzAE0EcwBhBHMAUwRzAFUCOQC5AjkAqgSsAHAErAByBKwAcARzAFoIHwBvBVb//QVWAJYFxwBmBccAngVWAKIE4wCoBjkAbQXHAKQCOQC/BAAANwVWAJYEcwCWBqoAmAXHAJwGOQBjBVYAngY5AFgFxwChBVYAXATjADAFxwChBVYACQeNABkFVgAJBVYABgTjACkCOQCLAjkAAAI5ACcDwQA2BHP/4QKqAFkEcwBKBHMAhgQAAFAEcwBGBHMASwI5ABMEcwBCBHMAhwHHAIgBx/+iBAAAiAHHAIMGqgCHBHMAhwRzAEQEcwCHBHMASAKqAIUEAAA/AjkAJARzAIMEAAAaBccABgQAAA8EAAAhBAAAKAKsADkCFAC8AqwALwSsAFcFVv/9BVb//QXHAGgFVgCiBccAnAY5AGMFxwChBHMASgRzAEoEcwBKBHMASgRzAEoEcwBKBAAAUARzAEsEcwBLBHMASwRzAEsCOQC9AjkAIwI5/+UCOQAJBHMAhwRzAEQEcwBEBHMARARzAEQEcwBEBHMAgwRzAIMEcwCDBHMAgwRzAEkDMwCABHMAawRzABsEcwBRAs0AbQRMAAEE4wCZBeUAAwXlAAMIAADhAqoA3gKqAD0EZABOCAAAAQY5AFMFtACaBGQATgRkAE0EZABNBHP//QScAKAD9AA4BbQAegaWAKEEZAAAAjEAAAL2AC8C7AAtBiUAfwcdAEQE4wCBBOMAngKqAOgErAByBGQAVARzAC4EZAAzBOUAGgRzAIYEcwCMCAAA7wVW//0FVv/9BjkAYwgAAIEHjQBSBHP//AgAAAACqgBTAqoARwHHAIABxwBsBGQATgP0AC8EAAAhBVYABgFW/jkEc//kAqoAXAKqAFwEAAAXBAAAFwRzAEkCOQC5AccAbAKqAEcIAAAlBVb//QVWAKIFVv/9BVYAogVWAKICOQCNAjn/4AI5AAQCOQAVBjkAYwY5AGMGOQBjBccAoQXHAKEFxwChAjkAxgKqABkCqgAGAqoAHQKqAC4CqgDlAqoAogKqAGsCqgA6AqoASwKqACgEcwAAAccAAwVWAFwEAAA/BOMAKQQAACgCFAC8Bcf//QRzAEkFVgAGBAAAIQVWAJ4EcwCHBKwAcgSsAKECqgBrAqoAGQKqACEGrABrBqwAawasACEEcwAABjkAbQRzAEICOQCxBVYAXAQAAD8FxwBmBAAAUAXHAGYEAABQBHMARgRr/+ECqgDuBVb//QRzAEoFVv/9BHMASgXHAJ4E6wBHBcf//QVWAKIEcwBLBVYAogRzAEsEcwCWAccAQgRzAJYCVQCIBHMAmgKsAIMFxwCcBHMAhwXHAJwEcwCHBjkAYwRzAEQFxwChAqoAhQXHAKECqgA8BVYAXAQAAD8E4wAwAjkAJATjADADAAAjBccAoQRzAIMFxwChBHMAgwTjACkEAAAoBOMAKQQAACgEaACkBjkAYAZiAFUEoABIBHQASAORAGIE8ABEAykALgUwAEgEa//hBAAAsALrAFIIwAAzCAAATwQAAJkIAABPBAAAmQgAAE8EAACYBAAAmAfVAWoFwACeBKsAcgTVAJ0ErABxBNUCIgTVAQUFq//pBQAByQWrAn4Fq//pBasCfgWr/+kFqwJ+Bav/6QWr/+kFq//pBav/6QWr/+kFqwHABasCfgWrAcAFqwHABav/6QWr/+kFq//pBasCfgWrAcAFqwHABav/6QWr/+kFq//pBasCfgWrAcAFqwHABav/6QWr/+kFq//pBav/6QWr/+kFq//pBav/6QWr/+kFq//pBav/6QWr/+kFq//pBav/6QWr/+kFq//pBav/6QWrAtYFqwBmBav/6gXV//8E1QCSCAAAAAfrATAH6wEgB+sBMAfrASAE1QCyBNUAgATVACoIKwGYCGsBuAdVABAGAAD0BgAAbwRAADoFQAA3BMAAPwQVAEAEAAAlBgAAVQXhAL8DjQCJBNX/2QGAAIAC1QCGBxUAYQKWAA8E1QCSAtYAgwLWAIME1QCyAtYAcAVW//0EcwBKBccAZgQAAFAFxwBmBAAAUAVWAKIEcwBLBVYAogRzAEsFVgCiBHMASwY5AG0EcwBCBjkAbQRzAEIGOQBtBHMAQgXHAKQEcwCHBccAHwRzAAYCOf/OAjn/zgI5/+QCOf/kAjn/9gI5//UCOQBLAccAGQQAADcBx/+iBVYAlgQAAIgEAACGBHMAlgHH//oFxwCcBHMAhwXJAKUEcwCLBjkAYwRzAEQGOQBjBHMARAXHAKECqgBrBVYAXAQAAD8E4wAwAjkADAXHAKEEcwCDBccAoQRzAIMFxwChBHMAgwXHAKEEcwCDB40AGQXHAAYFVgAGBAAAIQHHAIkFVv/9BHMASggAAAEHHQBEBjkAUwTjAIECOQC5B40AGQXHAAYHjQAZBccABgeNABkFxwAGBVYABgQAACEBxwCKAqr/4QRzABsEzQBaBqwAawasACIGrAAiBqwASgKqAOICqgBrAqoA3gKq/+oFV///Bkb/pwa0/6gDEv+oBjL/pwbY/6cGBf+nAcf/eAVW//0FVgCWBVj//gVWAKIE4wApBccApAI5AL8FVgCWBVgACwaqAJgFxwCcBTMAbQY5AGMFxwCkBVYAngTyAJQE4wAwBVYABgVWAAkGrwB/BfsAYQI5AAQFVgAGBKAASAORAGIEcwCLAccAawRgAIgEmgCMBAAAGQOHAEgEcwCLBHMAXAHHAIkEAACGBAAAGAScAKAEAAAaA5UAXARzAEQEjQCDA9sAVgRgAIgEMwARBbQAegY/AFcBx//JBGAAiARzAEgEYACIBj8AVwVXAKIG6wAyBFUAoQXAAGQFVgBcAjkAvwI5AAQEAAA3CHUADQgVAKQG1QAxBKkAoQUVAAoFwACgBVb//QVAAKcFVgCWBFUAoQVrAAAFVgCiB2MABwTVAE4FwAChBcAAoQSpAKEFQAASBqoAmAXHAKQGOQBjBcAAoAVWAJ4FxwBmBOMAMAUVAAoGFQBSBVYACQXrAJ8FVQBXB1UAoQeAAKEGVQAABxUAqAVAAKUFwABVCBUApAXHABoEcwBKBJUAWwRAAIgC6wCIBKsAAARzAEsFWv/7A6sAMgR4AIcEeACHA4AAhgSrABgFgACMBGsAiARzAEQEVQCIBHMAhwQAAFADqgAmBAAAIQaVAEsEAAAPBJUAigQrAEUGawCNBpUAjQUAACgFwACLBCsAhAQVADAGAACJBFUAHwRzAEsEcwAAAusAiQQVAEsEAAA/AccAiAI5AAkBx/+iB0AAEwaAAIMEcwAAA4AAhgQAACEEawCIA+kAoQNKAIgIAABBCJUAoAWFAC0AAAEBAAAAHgAAADEAAAAxAAABAQAAAH4AAAB+AAAAjAAAAIwAAAEBAAAAEAAAAQEAAAEhAxAAfQAAAIwCMwDSAAADCwAA/wQCOQC5BIEAaQRWADIDMQAZBBEALQTRAJYB+QCbAw8AXwTKAJsEuACMAfkAmwQTACgDsABQA7QAPATKAJsEzwBQAfkAmwLSADwEmABaBDwAGQSIAG4EXwBzA7EAGQPUAAoEZgCWBBMAKAWOAGQFJAAoA/IAmwPyAJsD8gCbAeMAWgNWAFoGhgCbAfn/rAQTACgEEwAoA7T/VwO0/1cESAAtBY4AZAWOAGQFjgBkBY4AZASBAGkEgQBpBIEAaQRWADIDMQAZBBEALQTRAJYCSwAAA0oAAAS4AIwCSwAABBMAKAOwAFADtAA8BM8AUALSADwEmABaBIgAbgRfAHMD1AAKBGYAlgQTACgFjgBkBSQAKAH5AJsEVgAyA7AAUARfAHMEmwA8AAD/3AAA/yUAAP/cAAD+UQKNAKsCjQCgAtoAQwNNAHkBqP+6AAAARgAAAEYAAABGAAAARgAAAEgAAABGAAAARgAAAEYENQF8BDUBLgQ1ALcENQCBBDUBLAQ1AL4ENQCvBDUAgQQ1AJoENQDbBDUAhQKNAMEENQCzBgABAAYAAQACQgA2BgABAAQ1AJ4ENQCYBDUAywYAAQAGAAEABgABAAYAAQAGAAEAAAAARgYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABRv/ugYAAQAGAAEABgABAAW1ADoFtQA6AfT/ugH0/7oGAAEABgABAAYAAQAGAAEABIEANgQ1ADYEPf+6BD3/ugPpAEoD6QBKBn8AFAd2ABQDJ/+6BB7/ugZ/ABQHdgAUAyf/ugQe/7oFGwAyBLUAJAMA//cGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAAAAAwAAAARgAAAEYAAABAAAAARgYAAQAGAAEAAAD/3AAA/lEAAP8WAAD/FgAA/xYAAP8WAAD/FgAA/xYAAP8WAAD/FgAA/xYAAP/cAAD/FgAA/9wAAP8gAAD/3ARzAEoIAAAABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAKNAH8CjQBdBgABAATuABUDTQB5AagADgHW/9wBqABWAdYAEAN1ADIDdQAyAagALQHWABMFGwAyBLUAJAH0/7oB9P+6AagAkwHWABMFtQA6BbUAOgH0/7oB9P+6AkIAAAMA//cFtQA6BbUAOgH0/7oB9P+6BbUAOgW1ADoB9P+6AfT/ugSBADYENQA2BD3/ugQ9/7oEgQA2BDUANgQ9/7oEPf+6BIEANgQ1ADYEPf+6BD3/ugKzAF8CswBfArMAXwKzAF8D6QBKA+kASgPpAEoD6QBKBpIAPgaSAD4EP/+6BD//ugaSAD4GkgA+BD//ugQ//7oIyQA+CMkAPgbF/7oGxf+6CMkAPgjJAD4Gxf+6BsX/ugSn/7oEp/+6BKf/ugSn/7oEp/+6BKf/ugSn/7oEp/+6BFoAKgOaADYENf+6Ayf/ugRaACoDmgA2BDX/ugMn/7oGTwAnBk8AJwIk/7oCGv+6BKcARgSnAEYCJP+6Ahr/ugTPAC0EzwAtAyf/ugMn/7oEDQBHBA0ARwGo/7oBqP+6ArQAIwK0ACMDJ/+6Ayf/ugQ1AEUENQBFAfT/ugH0/7oCQgA2AwD/9wOa/7oDJ/+6A3UAMgN1ADIFGwAyBLUAJAUbADIEtQAkAfT/ugH0/7oEWgBABM4ASQRaACYEzgA5BFoAUwTOAEoEWgBTBM4ASgYAAQAGAAEAAAAARgAAAEYGAAEABgABAAYAAQAAAABGAAAARgYAAQAGAAEAAAAASAAAAEYGAAEABgABAAYAAQAAAABGAAAARgAAAEYAAABGAAAAQAAAADAGAAEAAAAARgAAAEYGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQACjQDKAo0AxwKNAMYGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQABAP+6CAD/uhAA/7oG3ABjBT8ARAbVAKEFWwCDAAD93AAA/C8AAPymAAD+VAAA/NcAAP1zAAD+KQAA/g0AAP0RAAD8ZwAA/Z0AAPv1AAD8cgAA/tUAAP7VAAD/AgQbAKAGrABrBqwAGQAA/rYAAP1zAAD+CAAA/KYAAP5TAAD9EQAA+8gAAPr0AAD6rwAA/HIAAPuqAAD7agAA/PEAAPx9AAD73QAA/MEAAPuYAAD96gAA/oQAAP3CAAD88QAA/V8AAP52AAD+vAAA/OsAAP1sAAD9WAAA/JAAAP0VAAD8LAAA/BMAAPwSAAD7lgAA+5YBxwCIBVb//QRzAEoFVv/9BHMASgVW//0EcwBKBVb//QRzAEoFVv/9BHMASgVW//0EcwBKBVb//QRzAEoFVv/9BHMASgVW//0EcwBKBVb//QRzAEoFVv/9BHMASgVW//0EcwBKBVYAogRzAEsFVgCiBHMASwVWAKIEcwBLBVYAogRzAEsFVgCiBHMASwVWAKIEcwBLBVYAogRzAEsFVgCiBHMASwI5AGMBxwAfAjkAugHHAHwGOQBjBHMARAY5AGMEcwBEBjkAYwRzAEQGOQBjBHMARAY5AGMEcwBEBjkAYwRzAEQGOQBjBHMARAbcAGMFPwBEBtwAYwU/AEQG3ABjBT8ARAbcAGMFPwBEBtwAYwU/AEQFxwChBHMAgwXHAKEEcwCDBtUAoQVbAIMG1QChBVsAgwbVAKEFWwCDBtUAoQVbAIMG1QChBVsAgwVWAAYEAAAhBVYABgQAACEFVgAGBAAAIQVW//0EcwBKAjn/4gHH/7AGOQBjBHMARAXHAKEEcwCDBccAoQRzAIMFxwChBHMAgwXHAKEEcwCDBccAoQRzAIMAAP7+AAD+/gAA/v4AAP7+BFX//QLrAAwHYwAHBVr/+wSpAKEDgACGBKkAoQOAAIYFxwCkBGsAiARz//0EAAAUBHP//QQAABQFVgAJBAAADwVVAFcEKwBFBVUAoQRzAIcGBQBjBHMAVQY5AGAEcwBEBbUAOgH0/7oCJP+6Ahr/ugSnAEYB9ACeAfQAEAH0ABsB9AAQAfQAawH0//kCJ//OAAAADwAA//UCqgCkAqoApAAAAA4AAABWAAAAVgAA/88BqAAPAdb/vwGo//UB1v/NAagAHQHW//UBqACTAdYAEwN1ADIDdQAyA3UAMgN1ADIFGwAyBLUAJAW1ADoFtQA6AfT/ugH0/7oFtQA6BbUAOgH0/7oB9P+6BbUAOgW1ADoB9P+6AfT/ugW1ADoFtQA6AfT/ugH0/7oFtQA6BbUAOgH0/7oB9P+6BbUAOgW1ADoB9P+6AfT/ugW1ADoFtQA6AfT/ugH0/7oEgQA2BDUANgQ9/7oEPf+6BIEANgQ1ADYEPf+6BD3/ugSBADYENQA2BD3/ugQ9/7oEgQA2BDUANgQ9/7oEPf+6BIEANgQ1ADYEPf+6BD3/ugSBADYENQA2BD3/ugQ9/7oCswAyArMAMgKzAF8CswBfArMAXwKzAF8CswAyArMAMgKzAF8CswBfArMAXwKzAF8CswBfArMAXwKzADgCswA4ArMASQKzAEkD6QBKA+kASgPpAEoD6QBKA+kASgPpAEoD6QBKA+kASgPpAEoD6QBKA+kASgPpAEoD6QBKA+kASgPpAEoD6QBKBpIAPgaSAD4EP/+6BD//ugaSAD4GkgA+BD//ugQ//7oGkgA+BpIAPgQ//7oEP/+6CMkAPgjJAD4Gxf+6BsX/ugjJAD4IyQA+BsX/ugbF/7oEp/+6BKf/ugRaACoDmgA2BDX/ugMn/7oGTwAnBk8AJwZPACcCJP+6Ahr/ugZPACcGTwAnAiT/ugIa/7oGTwAnBk8AJwIk/7oCGv+6Bk8AJwZPACcCJP+6Ahr/ugZPACcGTwAnAiT/ugIa/7oEpwBGBKcARgSnAEYEpwBGCT4AMgk+ADIHQP+6B0D/ugZ/ABQHdgAUAyf/ugQe/7oEzwAtBM8ALQMn/7oDJ/+6BM8ALQTPAC0DJ/+6Ayf/ugTPAC0EzwAtAyf/ugMn/7oGfwAUB3YAFAMn/7oEHv+6Bn8AFAd2ABQDJ/+6BB7/ugZ/ABQHdgAUAyf/ugQe/7oGfwAUB3YAFAMn/7oEHv+6Bn8AFAd2ABQDJ/+6BB7/ugQNAEcEDQBHAaj/ugGo/7oEDQBHBA0ARwGo/7oBqP+6BA0ARwQNAEcBqP+6Aaj/ugQNAEcEDQBHAaj/ugGo/7oENQBFBDUARQH0/7oB9P+6BDUARQQ1AEUENQBFBDUARQQ1AEUENQBFAfT/ugH0/7oENQBFBDUARQSBADYENQA2BD3/ugQ9/7oCQgA2AwD/9wMaABoDGgAaAxoAGgN1ADIDdQAyA3UAMgN1ADIDdQAyA3UAMgN1ADIDdQAyA3UAMgN1ADIDdQAyA3UAMgN1ADIDdQAyA3UAMgN1ADIFG/+6BLX/ugUbADIEtQAkAfT/ugH0/7oDdQAyA3UAMgUbADIEtQAkAfT/ugH0/7oFGwAyBLUAJAZ/AEUGfwBFBn8ARQZ/AEUBqAAoAAD+KQAA/qIAAP8wAAD/HQAA/xIAAP+SAAD+fgj8ADIIrQAyAAD/tQAA/7YAAP7tAAD/ZAAA/n4AAP+fAY0AAAL2//0AAP6CAAD/EATNADIAAP9YAAD/WAAA/2QGkgA+BpIAPgQ//7oEP/+6CMkAPgjJAD4Gxf+6BsX/ugRaACoDmgA2BDX/ugMn/7oDTQB5ArQAIwJCADYB9P+6ApD/ugH0AC8B9AA7AfQAEgH0ALEB9ABtBn8AFAd2ABQB+QCbAAD+2QK8AAAD8gCbBFr/9QTO//UEWgBTBM4ASgRaAFMEzgBKBFoAUwTOAEoEWgBTBM4ASgRaAFMEzgBKBFoAUwTOAEoENQBxBDUArQRaAA8EzgAPBHMAFAYRABQFQACnBHMAhgVAAAoEcwAKBccAUQXHAGYEAABQBcf//QZ6ABQFQABKBHMARgR0AEgFVgBuBNUAUwTj/8QGOQBtBP4ADwcMAIcBxwCDAjkAHwVWAJYEAACIAccAFQQAABgHIACkBcf/uARzAIsGOQBgBvIAYwVXAEQGCQAUBHMAhgVWAJ4FVgBrBAAATwTyAJQDCwBEAjkAJATjABQCOQAkBOMAMAX7AGEFxwChBi4AEAQAACEE4wApBAAAKATjACkE4wAxBFwARARcAD8EcwA8BHMAVQOrADID5QAkBHMAhwIUALwDTgC8BKwAcgI5ALAKqgCeCccAnghkAEYIfwCWBqoAlgOcAIMJxwCcB44AnAYrAIcEcwBVBVb//QRzAEoAAP7+BVb//QRzAEoIAAABBx0ARAY5AG0EcwAaBjkAbQRzAEIFVgCWBAAAiAY5AGMEcwBEBjkAYwRzAEQE4wApBFwATAHH/6IKqgCeCccAnghkAEYGOQBtBHMAQghGAKQE8gCeBccAnARzAIcFVv/9BHMASgVW//0EcwBKBVYAogRzAEsFVgCiBHMASwI5/4oCOf9kAjkABAI5//YGOQBjBHMARAY5AGMEcwBEBccAoQKq/8wFxwChAqoAaAXHAKEEcwB2BccAoQRzAIMFVgBcBAAAPwTjADACOQAkBFwAUQN+ABMFxwCkBHMAhwWmAKQE1gBeBIYAXgTjACkEAAAoBVb//QRzAEoFVgCiBHMASwY5AGMEcwBEAAD+/QY5AGMEcwBEBjkAYwRzAEQGOQBjBHMARAVWAAYEAAAhBHMAVwRzAEgEcwCGBHMAhgQAABMEAABQBHMARgRzAEYEcwBVBekAVQOrAEkDqwAyBQ0AMgQPAEQCOf+5BHMAQgRzAEIEeABQBAIAGQTvABkEcwCLBHMAhwRzAIcBxwAZAccAVwLZAEQCngAAAm4AFAHHAIMEkwCDBqoAhAaqAIQGqgCHBHP/pgRzAIsEbACHBHMARAZTAEQGPwBXBGYARAKq/+QCqv/kAqr/5AKqAIUCqgCFAqoAhQKq/+QEVQCKBFUAigQAAD8Bx/+iAhT/uQHH/3ICywAAAjkADwI5ACQEcwAZBIwAVARgAIgEAAAaBccABgQAABgEKAAZBAAAKARUACgEXABMBFwAeQQAACQEAABQBAAAJAQAAFAGOQBjBEAAiAQPAEkEeABQBGsAiAMuAAAEAAAIAzsAiARzAEgEAAAkBAAAUAe3AEYHQABGCAsARgWzACQDbwAkBcAAJAYcABMFSgCDBQ8AgwPiAB4EOABjAxEAZAMRAGQBRv/OAesAZAHrAAAB6wAAAuoAZAPZAAACkQAAAYcAWgLXAF4BxwCAAccAbAHHAIoCqgD7AqoA+wLKADICygAyBKwAcASsAHAErABlBKwAZQKqASECqgDeAqoAWQKqASECqgAdAqoAWQKqAN4COQC2AjkAtgKqAPsCqgD7AqoApgKqAKYCqgCmAqoAHQKq/+ICqv/7ApQAAAFCAGQCuAAyAqAAAALKADIDEACWAxAAlgMQAJYDEACWAxAAlgKqAGICqgBiAqoAKAKqAB0CqgBHBFcAlgRXAJYEVwCWBFcAlgRXAEMEVwBDBFcAQwRXAEMEVwBDAxAAQwRXAC8EVwAvBFcALwRXAC8EVwAvAxAALwRXACUEVwAlBFcAJQRXACUEVwAlAxAALwRXABoEVwAaBFcAGgRXABoEVwAaAxAAGgRXAEIEVwBCBFcAQgRXAEIEVwBCAxAAQgRXAJYEVwCWBFcAlgRXAJYEVwBCBFcAQgRXAEIEVwBCBFcAQgMQAEIEVwAvBFcALwRXAC8EVwAvBFcALwMQAC8EVwAvBFcALwRXAC8EVwAvBFcALwMQAC8EVwAmBFcAJgRXACYEVwAmBFcAJgMQACYEVwBCBFcAQgRXAEIEVwBCBFcAQgMQAEIEVwCWBFcAlgRXAJYEVwCWBFcAQgRXAEIEVwBCBFcAQgRXAEIDEABCBFcAJgRXACYEVwAmBFcAJgRXACYDEAAmBFcAIwRXACMEVwAjBFcAIwRXACMDEAAjBFcALwRXAC8EVwAvBFcALwRXAC8DEAAvBFcASwRXAEsEVwBLBFcASwRXAEsDEABLBFcAlgRXAJYEVwCWBFcAlgRXAEIEVwBCBFcAQgRXAEIEVwBCAxAAQgRXABoEVwAaBFcAGgRXABoEVwAaAxAAGgRXACQEVwAkBFcAJARXACQEVwAkAxAAJARXAC8EVwAvBFcALwRXAC8EVwAvAxAALwRXAE4EVwBOBFcATgRXAE4EVwBOAxAATgRXAJYEVwCWBFcAlgRXAJYAAP7BAAD+xgAA/awAAP7YAAD/kgAA/ukAAP9MAAD+oAAA/sQAAP/OAAD/ZgAA/qAAAP7YAAD+2AAA/5cAAP+YAAD/mQAA//QAAP9CAAD/QgAA/0QAAP9fAAD+hwAA/+wAAP+mAAD/UQAA/1EAAP9RAAD+yQAA/xwAAAAAAAD+6QAA/0wAAP+TAAD/KgAA/1YAAP/OAAD+hwAA/rsAAP7EAAD+xAAA/tgAAP7YAAD+swAA/skAAP2tAAD+yAAA/rMAAP7JAAD9rQAA/hYAAP7mAAD/pgAA/ocAAP9EAAD+ugAA/yMAAP+aAAD9rAAA/ogAAAAAAAD+sAAA/5gAAP6TAAD/pgAA/ocAAP4cAAD/ZgAA/0QAAP6wAAD+sAAA/rAAAP8DAAD/UgAA/R8AAP9TAAD/UwAA/1MAAP61AAD+tQAA/8MAAP6uAAD+3AAA/scAAP7IAAD+3AAA/h4AAP9CAAD/UQAA/rcAAP6wAqoA3gKqAFkCqgD6BJoAcARgAAAGLgAUB6oAAAYuABQEewBMBj8AVwTPAEQGOQBjBHMARAXHAHAEAABQBOMAqAM7AIgE/wAABDwAMgYNAAoEnQBCByAApAaqAIQFZQBjBHMAiwVkAKQEAAAKBVYAawVWAGsE4AAFBMUAGQXlAF8EbgBEA7YAFANHACgEzwBEBJUAWwQAAFABx/+iBjkAYAOJAE0DiQBQBVYAogXAAKEEcwBLBHgAhwq0AG0E/gAQBjkAFATnABQHmQC/BbUAiAVYAAEEAAAGBy4AvwWQAIgGoQB4BXsAeghtAL8G8ACIBNUAZgOrAB8GXwA5BYIASAY5AGAEcwBEBm0ACQUMABoGbQAJBQwAGgiYAGMHLABEBqoAIATmABwJhwBtBtAAUAAA/jcKtABtBP4AEAXHAGYEAABQBAcAFAAA/qYAAP68AAD/mAAA/5gAAPwrAAD8TAXAAKEEeACHBUAABAQrABQFVgCeBHMAhwVdAKQEZACIBNUATgOrADIEqQAEA4AAAAXvACkESQAoBwkApAUvAIgJGACgBvYAiAYGAD4EKwAjBccAZgQAAFAE4wAwA6oAJgdnADEFhwAmBVUAVwQrAEUG5AAKBVQACgbkAAoFVAAKAjkAvwdjAAcFWv/7BVcAoQRoAIYFQAASBKsAGAXHAKQEawCIBccApARrAIgFVQBXBCsARQaqAJgFgACMAqoALgVW//0EcwBKBVb//QRzAEoIAAABBx0ARAVWAKIEcwBLBgUAYwRzAFUHYwAHBVr/+wTVAE4DqwAyBNUATgRcAEwFwAChBHgAhwXAAKEEeACHBjkAYwRzAEQGOQBgBHMARAXAAEoEFQArBRUACgQAACEFFQAKBAAAIQUVAAoEAAAhBVUAVwQrAEUHFQCoBcAAiwVAAEoEcwBGB78ASgcDAEYHpgBmBoYAUwVNAGYEEwBTB8MAEgdHABgIRgCkBwcAiAY5AG0EeABQBfkAMAVTACYAAP9DAAD+yQAA/3cAAP+wAAD/RwAA/1YAAP90AAD+1wAA/qwAAAAAAAD/UgAA/1YAAAAAAAD+rAAA/ZoAAAAAAAD/agAA/3wAAP9pAAD/VgAA/qwAAP9/AAD/VgAA/e8AAP9DAAD/aQAA/3wAAAAAAAD9rgAA/4wAAAECAAD+/gAA/v4AAP7fAAD+3wAA/1gAAP8gAAD+/gVW//0EcwBKBVYAlgRzAIYFVgCWBHMAhgVWAJYEcwCGBccAZgQAAFAFxwCeBHMARgXHAJ4EcwBGBccAngRzAEYFxwCeBHMARgXHAJ4EcwBGBVYAogRzAEsFVgCiBHMASwVWAKIEcwBLBVYAogRzAEsFVgCiBHMASwTjAKgCOQATBjkAbQRzAEIFxwCkBHMAhwXHAKQEcwCHBccApARzAIcFxwCTBHMAaAXHAKQEcwCHAjn/3wHH/5ICOQAgAjkABgVWAJYEAACIBVYAlgQAAIgFVgCWBAAAiARzAJYBxwB+BHMAlgHH/7kEcwCWAcf/pQRzAJYBx/+jBqoAmAaqAIcGqgCYBqoAhwaqAJgGqgCHBccAnARzAIcFxwCcBHMAhwXHAJwEcwCHBccAnARzAIcGOQBjBHMARAY5AGMEcwBEBjkAYwRzAEQGOQBjBHMARAVWAJ4EcwCHBVYAngRzAIcFxwChAqoAhQXHAKECqgCFBccAoQKqAF4FxwChAqoAJgVWAFwEAAA/BVYAXAQAAD8FVgBcBAAAPwVWAFwEAAA/BVYAXAQAAD8E4wAwAjkAJATjADACOQAkBOMAMAI5//8E4wAwAjkADgXHAKEEcwCDBccAoQRzAIMFxwChBHMAgwXHAKEEcwCDBccAoQRzAIMFVgAJBAAAGgVWAAkEAAAaB40AGQXHAAYHjQAZBccABgVWAAkEAAAPBVYACQQAAA8FVgAGBAAAIQTjACkEAAAoBOMAKQQAACgE4wApBAAAKARzAIcCOQADBccABgQAACEEcwBKAccAiQSgAEgEoABIBKAASASgAEgEoABIBKAASASgAEgEoABIBVb//QVW//0GggATBoIAEwaCABMGggATBoIAVgaCAFYDkQBiA5EAYgORAGIDkQBiA5EAYgORAGIGHgAABh4AAAdsAAAHbAAAB2wAAAdsAAAEcwCLBHMAiwRzAIsEcwCLBHMAiwRzAIsEcwCLBHMAiwaPAAAGjwAACB8AAAgfAAAIHwAACB8AAAgf//MIH//zAccAgQHHAIEBx/+bAcf/mwHH/+sBx//rAcf/ogHH/6IDAQAAAwEAAASRAAAEkQAABJEAAASRAAAEkf/zBJH/8wRzAEQEcwBEBHMARARzAEQEcwBEBHMARAadAAAGnQAACC0AAAgtAAAHyQAAB8kAAARgAIgEYACIBGAAiARgAIgEYACIBGAAiARgAIgEYACIBoIAAAeuAAAIEgAAB64ABgY/AFcGPwBXBj8AVwY/AFcGPwBXBj8AVwY/AFcGPwBXBl8AAAZfAAAH7wAAB+8AAAeLAAAHiwAAB4v//weL//8EoABIBKAASAORAGIDkQBiBHMAiwRzAIsBx//mAccAaARzAEQEcwBEBGAAiARgAIgGPwBXBj8AVwSgAEgEoABIBKAASASgAEgEoABIBKAASASgAEgEoABIBVb//QVW//0GggATBoIAEwaCABMGggATBoIAVgaCAFYEcwCLBHMAiwRzAIsEcwCLBHMAiwRzAIsEcwCLBHMAiwaPAAAGjwAACB8AAAgfAAAIHwAACB8AAAgf//MIH//zBj8AVwY/AFcGPwBXBj8AVwY/AFcGPwBXBj8AVwY/AFcGXwAABl8AAAfvAAAH7wAAB4sAAAeLAAAHi///B4v//wSgAEgEoABIBKAASASgAEgEoABIBKAASASgAEgFVv/9BVb//QVW//0FVv/9BVb//QKqAOUCqgD9AqoA5QKqAAYCqgAGBHMAiwRzAIsEcwCLBHMAiwRzAIsGggAABoIAAAbzAAAG8wAABccApAKqABMCqgATAqoABgHH/7sBx/+rAcf/ygHH/8oBx/+TAcf/kwI5ABoCOf/1A2UAAANlAAACqgATAqoAEwKqAAYEYACIBGAAiARgAIgEYACIBI0AgwSNAIMEYACIBGAAiAVWAAYFVgAGBuYAAAcYAAAGHgAAAqr/6gKq/+oCqgBZBj8AVwY/AFcGPwBXBj8AVwY/AFcHZQAABp0AAAcnAAAGXwAABfsAYQKqAN4CqgDlBHMADQXHAGYFxwBmBqoAhwXHACQJUAChB40AGQVWAB8E4wAwCAAAKQQAADAEwQBmAAD/UwAA/1MAAP9TAAD/UwHHABkBx/+iBCsABQVWABEFdABGAsv/owV6AIcC8P/IBX8ACgV/AAoCqgCEAqoAhAKqAMkCqgDJAqoAoAKqAFkCqv+vAqoAOgKqAAYCOQC5AqoAqQKqAKkCqgCpAqoAqQMuAB4DLgAeAqoAOgAA/3MAAP+lAAD+2AAA/yMAAP9yAAD/cgAA/ucAAP+lAAD/UwAA/1MAAP9TBVYAngRzAIcD+AAZBfsAGQcdAEQEQAAZBAAAUARpAIcEaQAZA+sAhwOrADIBxwCIA2EAQQQAAIgDNgAQBYAAjAR4AIcEcwBEBAAAEwTeAEQE3gBEBN4ADQeNAFADqABEBHMARARzAEQEKwCEBFUAHwRVAB8DqgAmBGAAiATGAEQF3gBEBMYARAQAABoFxwAGBAAAKAOrADIDawA/BNsAHwLrAIgEAAAaBFUAiAQrAIQFtAB6BKsAGAOgAAAFTwAAA1EAMgNR/9EDmAAyA0gAMgNIADID+AAyA24AMgFWAGkChAAtA2YAMgLQADIEFQAyA3EAMgNvADIEGAAyAw8AMgNZADIDnAAyA3YAMQNvADIE+wAAAvoAMgL6ADIDBAAyBMwAMgMFAGQDBQAyAvkAMgL5ADICjAAyAowAMgMEADIBQgBkArYAZASVAGQDDwBkAwUAMgLVADIDBQAyAwUAMgMGAGQBwgAyAw8AZANCADIElQBkApIAAAMgAAADFQBkApIAAAMGADIDhQAyAr8AAAFCAGQB6wBkAw8AZAKSAAADFQBkApIAAAMJADIDhQAyAr8AAAXtAEYKZgBGBhMARgaJ/7oFQf+6AekAPARaABEAAP8NAAD/NQAA/s4AAP63AAD+yQAA/88AAP9PAAD/ngAA/soCswBfArMAXwPpAEoD6QBKA5r/ugMn/7oDmv+6Ayf/ugWtAGkFPQAtBf0AlgTcAFAE4AA8BfYAmwU/ACgGUAAoBKwAcgAA/jsAAP5mAAD+ZgRz//wCqgBTAtX/zgGo/7oBqP+6Aaj/ugGo/7oGWAAVCcUARwQAAAAIAAAABAAAAAgAAAACqwAAAgAAAAFVAAAEcwAAAjkAAAGaAAAAqwAAAAAAAAXlAAMFxwBmBqoAmAWAAIwHRACDBxgARgcYAEgFVv/9BccAZgQAABQEcwAKBOMAMAQAAE8EAAAoBKUAHQAAAQIAAP9CAAD+vwAA/zoAAP9TBI0ACgXHAFEFxwBmBccAUQRVAKEC6wCIAAD/QwAA/wQAAP+sAtIAlgAA/zcCGv+6AlAAHgAA/zoAAP9bAAD/XwAA/34AAP+UAAD/SgAA/pwFtQA6BbUAOgH0/5YB9P+WBbUAOgW1ADoB9P+6AfT/ugW1ADoFtQA6AfT/ugH0/7oFtQA6BbUAOgH0/7oB9P+6BbUAOgW1ADoB9P+6AfT/ugW1ADoFtQA6AfT/ugH0/7oFtQA6BbUAOgH0/7oB9P+6BIEANgQ1ADYEPf+6BD3/ugSBADYENQA2BD3/ugQ9/7oCswAyArMAMgKzAF8CswBfA+kASgPpAEoGkgA+BpIAPgQ//7oEP/+6BFoAKgOaADYENf+6Ayf/ugRaACoDmgA2BDX/ugMn/7oEWgAqA5oANgQ1/7oDJ/+6Bk8AJwZPACcCJP+6Ahr/ugZPACcGTwAnAiT/ugIa/7oGfwAUB3YAFAMn/7oEHv+6Bn8AFAd2ABQDJ/+6BB7/ugZ/ABQHdgAUAyf/ugQe/7oCtAAjArQAIwMn/7oDJ/+6ArQAIwK0ACMDJ/+6Ayf/ugQ1AEUENQBFAfT/ugH0/7oENQBFBDUARQH0/7oB9P+6BDUARQQ1AEUB9P+6AfT/ugQNAEcEDQBHAaj/ugGo/7oD6QBKA+kASgPpAEoD6QBKBpIAPgaSAD4EP/+6BD//ugRz/5MEcwBGAjn/vwaq/9UEc/+3BHP/kQKq/6QCqv+kBAD//wI5/7kEAAAoBHMAiQMLAGQEdABIBkkAJAHHABkBxwAZBHMAHgRgAB4EjAAKBHMAhgRzAEYCOQATBbQAQgQAAIgBx//8BqoAhwRzAIsEcwCHAqr/+wQAAD8DGP+iBAAAGgQAAA8EAAAoBHMASgRzAEgEcwBGBHMASwOrAEkDqwAyBTQAVQHHAIgEAAATAcf/ogRzAIMEXABMAwQAZALVADICyQAzAvwAMgKMADIB1QAyAdUAAAMEADIDEQBkAUIAGQFCAGQBQgBkAUIAGQIqAAABQgBkAUIACQIzAGQEkwBkBJMAZAMP/8kDDwBkAw4AZAMFADIDAAAyArgAMgFC/8oBwgAyAw8AHQMaADIDBgBkAtQAZAKSAAAC3gAyAt4AMgLeADIC9AAyAuoAMgAA/rwAAP68AAD/cwAA/qkCOQC5AvoAMgL5ADIDBQAyAqAAAAL5ADIGOQBtBVb//QRzAA8FxwBmAqoAQQSgAEgEoABIBKAASASgAEgEoABIBKAASASgAEgEoABIAcf/mwHH/6sBx/+bAcf/qwHH/5sBx/+7Acf/mwHH/7sEYACIBGAAiARgAIgEYACIBGAAiARgAIgEYACIBGAAiAHH/6sBx/+rAcf/uwHH/7sEYACIBGAAiARgAIgEYACIBFoAUwTOAEoDoAATBVYAEQXHACkFWAALBVYAogRzAEsEAAAzAcf/ogXmAGMEcwBIBccAAAKqAA8FVgAGBAAAIQQAABMEAABQBAAAEwHHAIMEVf/9AusAAQVWAAkEAAAPBVYACQQAAA8E1QBTA6sASQVAABIEqwAYAAD+xgAA/tQAAP7GAAD+1AAA/l8AAP5fAAD/cgAA/3MAAP7nB4sACgPrAEwEAAATBHMACgHHABUEc//0BVYAEQXHAKEEcwAZAjn/iwXHAKQEcwCHBVYAlgQAAIgE4wApBAAAKAQAADsEngCkA2cAiAUwAEgAAP9TAAD/vAAA/v4AAP7+AAD+pAAA/qQBxwCIBckApQXHAJwFyQClAAD+zQAA/0gAAP7JAAD+zgAA/sUAAP7QAAD+0QAA/u4AAP7WAAD+3AAA/dkGOQBYBHMASAeNABkFxwAGBZ8ApAAA/rkF3ABjBMYACQhMABkGugAGAjkAuQOAAHIBhwBaAYcAWgQAAJkEAACZAjkAsAI5ALACOQCwAqoAGQTjADAEcwBQBHMADwRzABwGWwCHBkoATAAAAAAAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAAAYgAAAGIAAABiAAEAAA1dAPIAPACdAAcAAgAQAC8AVgAABKz//wAFAAIAAAAUAPYAAQAAAAAAAAAQAAAAAQAAAAAAAQAMABAAAQAAAAAAAgAHABwAAQAAAAAAAwAIACMAAQAAAAAABAAMACsAAQAAAAAABQAMADcAAQAAAAAABgAAAEMAAQAAAAAABwAHAEMAAQAAAAAACAAHAEoAAQAAAAAACQAHAFEAAwABBAkAAAAgAFgAAwABBAkAAQAYAHgAAwABBAkAAgAOAJAAAwABBAkAAwAQAJ4AAwABBAkABAAYAK4AAwABBAkABQAYAMYAAwABBAkABgAAAN4AAwABBAkABwAOAN4AAwABBAkACAAOAOwAAwABBAkACQAOAPpPcmlnaW5hbCBsaWNlbmNlQk9HQUhQK0FyaWFsVW5rbm93bnVuaXF1ZUlEQk9HQUhQK0FyaWFsVmVyc2lvbiAwLjExVW5rbm93blVua25vd25Vbmtub3duAE8AcgBpAGcAaQBuAGEAbAAgAGwAaQBjAGUAbgBjAGUAQgBPAEcAQQBIAFAAKwBBAHIAaQBhAGwAVQBuAGsAbgBvAHcAbgB1AG4AaQBxAHUAZQBJAEQAQgBPAEcAQQBIAFAAKwBBAHIAaQBhAGwAVgBlAHIAcwBpAG8AbgAgADAALgAxADEAVQBuAGsAbgBvAHcAbgBVAG4AawBuAG8AdwBuAFUAbgBrAG4AbwB3AG4AAAADAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAuQBUAyizJhgf0LwDKQDgAykAAgMpsisdH7kDJwMdsjsfQLgDI7MSFTIPQS0DIAABAC8DIAABACADIABvAyAArwMgAL8DIAAEAF8DHgABABADHgB/Ax4AgAMeAK8DHgC/Ax4A0AMeAAYAAAMeABADHgAgAx4AbwMeAJ8DHgDgAx4ABgMdAxyyIB8QQScDGQB/AxkAAgAPAxcA7wMXAP8DFwADAB8DFwAvAxcATwMXAF8DFwCPAxcAnwMXAAYADwMXAF8DFwBvAxcAfwMXAL8DFwDwAxcABgBAAxeykjNAuAMXsoszQLgDF7NqbDJAuAMXsmEzQLgDF7NcXTJAuAMXs1dZMkC4AxezTVEyQLgDF7NESTJAuAMXsjozQLgDF7MxNDJAuAMXsy5CMkC4AxezJywyQLgDF7MSJTKAuAMXswoNMsBBFgMWANADFgACAHADFgABAsQADwEBAB8AoAMVALADFQACAwYADwEBAB8AQAMSsyQmMp+/AwQAAQMCAwEAZAAf/8ADAbINETJBCgL/Au8AEgAfAu4C7QBkAB//wALtsw4RMp9BSgLiAK8C4gC/AuIAAwLiAuIC4QLhAH8C4AABABAC4AA/AuAAnwLgAL8C4ADPAuAA7wLgAAYC4ALgAt8C3wLeAt4ADwLdAC8C3QA/At0AXwLdAJ8C3QC/At0A7wLdAAcC3QLdABAC3AABAAAC3AABABAC3AA/AtwAAgLcAtwAEALbAAEC2wLbAA8C2gABAtoC2v/AAtOyNzkyuf/AAtOyKy8yuf/AAtOyHyUyuf/AAtOyFxsyuf/AAtOyEhYyuALSsvkpH7kDJgMcsjsfQLsDIgA+ADMDIrIlMR+4AxiyPGkfuALjsyArH6BBMALUALAC1AACAAAC1AAQAtQAIALUAFAC1ABgAtQAcALUAAYAYALWAHAC1gCAAtYAkALWAKAC1gCwAtYABgAAAtYAEALWACACygAgAswAIALWADAC1gBAAtYAUALWAAgC0LIgKx+4As+yJkIfQRYCzgLHABcAHwLNAsgAFwAfAswCxgAXAB8CywLFABcAHwLJAsUAHgAfAsoCxrIeHwBBCwLGAAACxwAQAsYAEALHAC8CxQAFAsGzJBIf/0ERAr8AAQAfAr8ALwK/AD8CvwBPAr8AXwK/AI8CvwAGAr8CIrJkHxJBCwK7AMoIAAAfArIA6QgAAB8CpgCiCABAah9AJkNJMkAgQ0kyQCY6PTJAIDo9Mp8gnyYCQCaWmTJAIJaZMkAmjpIyQCCOkjJAJoSMMkAghIwyQCZ6gTJAIHqBMkAmbHYyQCBsdjJAJmRqMkAgZGoyQCZaXzJAIFpfMkAmT1QyQCBPVDK4Ap63JCcfN09rASBBDwJ3ADACdwBAAncAUAJ3AAQCdwJ3AncA+QQAAB8Cm7IqKh+4AppAKykqH4C6AYC8AYBSAYCiAYBlAYB+AYCBAYA8AYBeAYArAYAcAYAeAYBAAYC7ATgAAQCAAUC0AYBAAYC7ATgAAQCAATlAGAGAygGArQGAcwGAJgGAJQGAJAGAIAE3QLgCIbJJM0C4AiGyRTNAuAIhs0FCMkC4AiGzPT4yD0EPAiEAPwIhAH8CIQADAL8CIQDPAiEA/wIhAAMAQAIhsyAiMkC4AiGzGR4yQLgCIrMqPzJAuAIhsy46Mm9BSALDAH8CwwCPAsMA3wLDAAQALwLDAGACwwDPAsMAAwAPAsMAPwLDAF8CwwDAAsMA7wLDAP8CwwAGAN8CIgABAI8CIgABAA8CIgAvAiIAPwIiAF8CIgB/AiIA7wIiAAYAvwIhAO8CIQACAG8CIQB/AiEArwIhAAMALwIhAD8CIQBPAiEAAwLDAsMCIgIiAiECIUAdEBwQKxBIA48cAQ8eAU8e/x4CNwAWFgAAABIRCBG4AQ229w349w0ACUEJAo4CjwAdAB8CkAKPAB0AHwKPsvkdH7gBmLImux9BFQGXAB4EAQAfATkAJgElAB8BOABzBAEAHwE1ABwIAQAfATQAHAKrAB8BMrIcVh+4AQ+yJiwfugEOAB4EAbYf+RzkH+kcuAIBth/oHLsf1yC4BAGyH9UcuAKrth/UHIkfyS+4CAGyH7wmuAEBsh+6ILgCAbYfuRw4H63KuAQBsh+BJrgBmrIffia4AZq2H30cRx9rHLgEAbIfZSa4AZqyH15zuAQBQA8fUiZaH0gciR9EHGIfQHO4CAG2Hz8cXh88JrgBmrIfNRy4BAG2HzAcux8rHLgEAbYfKhxWHykcuAEBsh8jHrgEAbIfVTe4AWhALAeWB1gHTwc2BzIHLAchBx8HHQcbBxQIEggQCA4IDAgKCAgIBggECAIIAAgUuP/gQCsAAAEAFAYQAAABAAYEAAABAAQQAAABABACAAABAAIAAAABAAACAQgCAEoAsBMDSwJLU0IBS7DAYwBLYiCw9lMjuAEKUVqwBSNCAbASSwBLVEKwOCtLuAf/UrA3K0uwB1BbWLEBAY5ZsDgrsAKIuAEAVFi4Af+xAQGOhRuwEkNYuQABARGFjRu5AAEBKIWNWVkAGBZ2Pxg/Ej4ROUZEPhE5RkQ+ETlGRD4ROUZEPhE5RmBEPhE5RmBEKysrKysrKysrKysYKysrKysrKysrKysYKx2wlktTWLCqHVmwMktTWLD/HVlLsJNTIFxYuQHyAfBFRLkB8QHwRURZWLkDPgHyRVJYuQHyAz5EWVlLuAFWUyBcWLkAIAHxRUS5ACYB8UVEWVi5CB4AIEVSWLkAIAgeRFlZS7gBmlMgXFi5ACUB8kVEuQAkAfJFRFlYuQkJACVFUli5ACUJCURZWUu4BAFTIFxYsXMkRUSxJCRFRFlYuRcgAHNFUli5AHMXIERZWUu4BAFTIFxYscolRUSxJSVFRFlYuRaAAMpFUli5AMoWgERZWUuwPlMgXFixHBxFRLEeHEVEWVi5ARoAHEVSWLkAHAEaRFlZS7BWUyBcWLEcHEVEsS8cRURZWLkBiQAcRVJYuQAcAYlEWVlLuAMBUyBcWLEcHEVEsRwcRURZWLkN4AAcRVJYuQAcDeBEWVkrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrK2VCKysBsztZY1xFZSNFYCNFZWAjRWCwi3ZoGLCAYiAgsWNZRWUjRSCwAyZgYmNoILADJmFlsFkjZUSwYyNEILE7XEVlI0UgsAMmYGJjaCCwAyZhZbBcI2VEsDsjRLEAXEVUWLFcQGVEsjtAO0UjYURZs0dQNDdFZSNFYCNFZWAjRWCwiXZoGLCAYiAgsTRQRWUjRSCwAyZgYmNoILADJmFlsFAjZUSwNCNEILFHN0VlI0UgsAMmYGJjaCCwAyZhZbA3I2VEsEcjRLEAN0VUWLE3QGVEskdAR0UjYURZAEtTQgFLUFixCABCWUNcWLEIAEJZswILChJDWGAbIVlCFhBwPrASQ1i5OyEYfhu6BAABqAALK1mwDCNCsA0jQrASQ1i5LUEtQRu6BAAEAAALK1mwDiNCsA8jQrASQ1i5GH47IRu6AagEAAALK1mwECNCsBEjQgArdHVzdQAYRWlERWlERWlEc3Nzc3R1c3R1KysrK3R1KysrKytzc3Nzc3Nzc3Nzc3Nzc3Nzc3Nzc3Nzc3NzKysrRbBAYURzdAAAS7AqU0uwP1FaWLEHB0WwQGBEWQBLsDpTS7A/UVpYsQsLRbj/wGBEWQBLsC5TS7A6UVpYsQMDRbBAYERZAEuwLlNLsDxRWlixCQlFuP/AYERZKysrKysrKysrKysrKysrKysrdSsrKysrKytDXFi5AIACu7MBQB4BdABzWQOwHktUArASS1RasBJDXFpYugCfAiIAAQBzWQArdHMBKwFzKysrKysrKytzc3NzKysrKysAKysrKysrAEVpRHNFaURzRWlEc3R1RWlEc0VpREVpREVpRHN0RWlERWlEcysrKysrcysAK3MrdHUrKysrKysrKysrKysrK3N0dXMrc3R1c3R1KysrdCsrAAA=); }&#xA;</svg:style><svg:clipPath id="clippath4" transform=""><svg:path d="M 200.22 566.48 L 394.978 566.48 L 394.978 754.036 L 200.22 754.036 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="none" clip-rule="nonzero"></svg:path></svg:clipPath><svg:clipPath id="clippath5" transform=""><svg:path d="M 200.22 566.48 L 394.978 566.48 L 394.978 754.036 L 200.22 754.036 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="none" clip-rule="nonzero"></svg:path></svg:clipPath></svg:defs><svg:g transform=""><svg:text transform="matrix(10.9755 0 0 10.98 294.66 795.7403) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_3" font-size="1px" y="0"></svg:tspan><svg:tspan x="0" y="0" font-family="g_font_3" font-size="1px" fill="rgb(0,0,0)">5</svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="0" x="0.5576" fill="rgb(0,0,0)"> </svg:tspan></svg:text><svg:text transform="matrix(7.9767 0 0 7.98 49.62 38.6603) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_2" font-size="1px" y="0" x="0 0.7375 1.016 1.7385 2.461 3.0175 3.685 4.3525 4.631 5.1875 5.744 6.308 6.872 27.5574 28.1139 28.6704 29.2269 29.7834 30.0619 30.6184 31.1749 31.4609 32.2394 32.5179 33.2404 33.5189 34.0754 34.6394" fill="rgb(0,0,0)">© UCLES 2017 0439/11/O/N/17 </svg:tspan></svg:text><svg:text transform="matrix(10.9755 0 0 10.98 491.28 38.6603) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_3" font-size="1px" y="0" x="0 0.3341 0.9462 1.5583 1.9484 2.5605 2.8395 3.4516 4.0087 4.5658" fill="rgb(0,0,0)">[Turn over</svg:tspan></svg:text><svg:text transform="matrix(7.9767 0 0 7.98 545.7 38.6603) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_2" font-size="1px" y="0" x="0" fill="rgb(0,0,0)"> </svg:tspan></svg:text><svg:text transform="matrix(10.9755 0 0 10.98 49.62 769.4603) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_3" font-size="1px" y="0" x="0 0.5575" fill="rgb(0,0,0)">10</svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="0" x="1.1152 1.9354 2.6038 2.8272 3.3846 3.886 4.1654 4.4998 4.7232 5.2246 5.448 5.7274 6.2288 6.5078 6.7312 7.2326 7.5061 8.0635 8.6209 9.1223 9.6237 10.1811 10.7385 11.0175 11.2969 11.8543 12.1887 12.7407 13.2981 13.8555 14.4129 14.6919 15.1933 15.7507 16.3081 16.8095 17.3669 17.9243 18.1978 18.5313 19.0887 19.3681 19.9255 20.4829 20.7619 21.3193 21.8767 22.4341 22.9915 23.5489 24.1063 24.6077 24.8867 25.3881 25.9455 26.5029 26.7263 27.2837 28.1181 28.3971 28.8985 29.4559 29.6793 30.2367 30.5711 30.7945 31.3519 31.9093 32.1887 32.4677 32.7471 33.3045 33.8619 34.1963 34.4698 34.7488 35.3062 35.5296 36.087 36.5884 36.8678 37.2022 37.7596 38.317 38.8744 39.3758 39.6493 40.2067 40.5411 41.0985 41.3775 41.9349 42.4363 42.9937 43.5511 43.8246" fill="rgb(0,0,0)"> Electricity is passed through concentrated aqueous sodium chloride. Inert electrodes are used. </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="1.153" x="0" fill="rgb(0,0,0)"> </svg:tspan></svg:text></svg:g><svg:g transform=""><svg:path d="M 200.22 566.48 L 394.978 566.48 L 394.978 754.036 L 200.22 754.036 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="none" clip-rule="nonzero"></svg:path></svg:g><svg:g clip-path="url(#clippath4)"><svg:g transform=""><svg:path d="M 200.22 566.48 L 394.978 566.48 L 394.978 754.036 L 200.22 754.036 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="none" clip-rule="nonzero"></svg:path></svg:g><svg:g transform=""><svg:path d="M 220.19 673.229 L 202.367 673.229 L 201.857 608.464 C 227.828 570.543 203.385 579.706 227.828 570.543 C 264.747 570.543 248.452 562.908 264.747 570.543 C 290.718 602.609 285.88 579.197 290.718 602.609 L 291.004 673.229 L 273.182 673.229 L 272.385 652.613 L 272.131 605.664 C 246.924 585.304 269.076 585.304 246.924 585.304 C 220.19 608.464 222.481 584.541 220.19 608.464 L 220.19 673.229" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(226,226,227)"></svg:path><svg:path d="M 272.661 688.372 L 272.661 610.266 C 272.661 603.6 270.063 597.329 265.346 592.615 C 260.629 587.901 254.359 585.304 247.688 585.304 L 245.182 585.304 C 238.511 585.304 232.241 587.901 227.525 592.615 C 222.807 597.329 220.21 603.6 220.21 610.266 L 220.21 688.372 C 221.463 690.662 219.808 690.026 221.463 690.662 M 290.992 688.372 L 290.992 610.266 C 290.992 586.361 271.604 566.98 247.688 566.98 L 245.182 566.98 C 221.266 566.98 201.878 586.361 201.878 610.266 L 201.878 688.372 C 200.457 690.917 202.111 690.026 200.457 690.917 M 290.974 688.372 C 292.226 690.662 290.571 690.026 292.226 690.662 M 272.641 688.372 C 271.22 690.917 272.875 690.026 271.22 690.917" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.999px" stroke-dasharray="" stroke-dashoffset="0px" fill="none" stroke="rgb(43,46,52)"></svg:path></svg:g></svg:g><svg:g transform=""><svg:path d="M 208.986 706.824 L 213.569 706.824 L 213.569 644.725 L 208.986 644.725 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(43,46,52)"></svg:path><svg:path d="M 208.986 644.725 L 213.569 644.725 L 213.569 706.824 L 208.986 706.824 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.999px" stroke-dasharray="" stroke-dashoffset="0px" fill="none" stroke="rgb(43,46,52)"></svg:path><svg:path d="M 279.26 706.824 L 283.843 706.824 L 283.843 644.725 L 279.26 644.725 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.999px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(43,46,52)"></svg:path><svg:path d="M 279.26 644.725 L 283.843 644.725 L 283.843 706.824 L 279.26 706.824 Z M 248.218 739.909 L 281.691 739.909 L 281.691 704.31 M 211.283 705.805 L 211.283 739.909 L 245.386 739.909" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.999px" stroke-dasharray="" stroke-dashoffset="0px" fill="none" stroke="rgb(43,46,52)"></svg:path><svg:path d="M 220.19 674.319 C 220.19 673.111 217.411 673.229 217.411 673.229 L 204.656 673.229 C 201.878 674.319 201.878 673.111 201.878 674.319 M 290.955 674.319 C 290.955 673.111 288.176 673.229 288.176 673.229 L 275.421 673.229 C 272.643 674.319 272.643 673.111 272.643 674.319" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="none" stroke="rgb(43,46,52)"></svg:path><svg:text transform="matrix(10.9966 0 0 10.9918 200.6037 709.0696) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_6" font-size="1px" y="0" x="0 7.7565" fill="rgb(43,46,52)">+–</svg:tspan><svg:tspan font-family="g_font_6" font-size="1px" y="7.5076" x="10.3376 10.8376 11.3936 11.9496 12.4496 13.0056 13.5616 13.8396 14.1726 14.7286 15.0066 15.5626" fill="rgb(43,46,52)">concentrated</svg:tspan><svg:tspan font-family="g_font_6" font-size="1px" y="8.5985" x="10.3376 10.8936 11.4496 12.0056 12.5616 13.1176 13.6736 14.1736 14.4516 14.9516 15.5076 16.0636 16.2856 16.8416" fill="rgb(43,46,52)">aqueous sodium</svg:tspan><svg:tspan font-family="g_font_6" font-size="1px" y="9.6894" x="10.3376 10.8376 11.3936 11.6156 12.1716 12.5046 12.7266 13.2826" fill="rgb(43,46,52)">chloride</svg:tspan></svg:text></svg:g><svg:g transform=""><svg:path d="M 200.22 566.48 L 394.978 566.48 L 394.978 754.036 L 200.22 754.036 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="none" clip-rule="nonzero"></svg:path></svg:g><svg:g clip-path="url(#clippath5)"><svg:g transform=""><svg:path d="M 200.22 566.48 L 394.978 566.48 L 394.978 754.036 L 200.22 754.036 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="none" clip-rule="nonzero"></svg:path></svg:g><svg:g transform=""><svg:path d="M 282.123 620.656 L 311.283 629.129" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.5px" stroke-dasharray="" stroke-dashoffset="0px" fill="none" stroke="rgb(43,46,52)"></svg:path><svg:path d="M 245.312 725.71 L 245.312 754.037 M 248.145 732.792 L 248.145 746.954" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.999px" stroke-dasharray="" stroke-dashoffset="0px" fill="none" stroke="rgb(43,46,52)"></svg:path></svg:g></svg:g><svg:g transform=""><svg:text transform="matrix(10.9755 0 0 10.98 395.22 566.3604) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_2" font-size="1px" y="0"></svg:tspan><svg:tspan x="0" y="0" font-family="g_font_2" font-size="1px" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="0.929" x="-31.4882" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="2.0875" x="-29.553 -28.6078 -28.0506 -27.4934 -27.2142 -26.9352 -26.712 -26.2108 -25.9318 -25.6526 -25.0954 -24.7674 -23.9365 -23.3793 -22.8221 -22.5431 -21.9859 -21.7067 -21.4277 -21.1485 -20.5913 -20.0341 -19.7551 -19.1979 -18.6407 -18.0835 -17.5263 -17.2471 -17.0239 -16.5227 -15.9655 -15.6865 -15.1293 -14.9061 -14.3489 -13.8477 -13.5685 -13.2343 -12.6771 -12.1199 -11.5627 -11.0055" fill="rgb(0,0,0)">What is formed at the negative electrode? </svg:tspan><svg:tspan font-family="g_font_3" font-size="1px" y="4.235" x="-29.553 -28.8316" fill="rgb(0,0,0)">A </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="4.235" x="-27.6178 -27.1161 -26.5584 -26.3347 -25.777 -25.4423 -25.2186 -24.6609 -24.1089" fill="rgb(0,0,0)">chlorine </svg:tspan><svg:tspan font-family="g_font_3" font-size="1px" y="6.2077" x="-29.553 -28.8316" fill="rgb(0,0,0)">B </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="6.2077" x="-27.6178 -27.0609 -26.56 -26.0031 -25.6692 -25.1123 -24.5554 -23.9985 -23.4416" fill="rgb(0,0,0)">hydrogen </svg:tspan><svg:tspan font-family="g_font_3" font-size="1px" y="8.1804" x="-29.553 -28.8316" fill="rgb(0,0,0)">C </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="8.1804" x="-27.6178 -27.0616 -26.5614 -26.0612 -25.505 -24.9488 -24.3859" fill="rgb(0,0,0)">oxygen </svg:tspan><svg:tspan font-family="g_font_3" font-size="1px" y="10.1531" x="-29.553 -28.8316" fill="rgb(0,0,0)">D </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="10.1531" x="-27.6178 -27.1166 -26.5594 -26.0022 -25.779 -25.2218 -24.3876" fill="rgb(0,0,0)">sodium </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="11.3006" x="-31.4882" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="12.4536" x="-31.4882" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_3" font-size="1px" y="13.6066" x="-31.4882 -30.9307" fill="rgb(0,0,0)">11</svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="13.6066" x="-30.373 -29.5528 -28.9406 -28.2174 -27.6602 -27.3812 -26.88 -26.3228 -25.7656 -24.9314 -24.7082 -24.207 -23.6498 -23.4266 -23.1476 -22.5904 -22.2562 -21.699 -21.1978 -20.6406 -20.1394 -19.6382 -19.0862 -18.585 -18.306 -17.7488 -17.4146 -16.8574 -16.5784 -16.0212 -15.464 -14.9628 -14.4616 -14.1274 -13.9042 -13.347 -12.7898 -12.2326 -11.9534" fill="rgb(0,0,0)"> Two chemical processes are described. </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="14.7596" x="-31.4882" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_9" font-size="1px" y="15.9126" x="-25.6771" fill="rgb(0,0,0)">●</svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="15.9126" x="-25.0703 -23.7363 -23.0132 -22.4561 -22.122 -21.8989 -21.3418 -20.7847 -20.5057 -20.2266 -19.6695 -19.1124 -18.8334 -18.3323 -17.7752 -16.9411 -16.384 -15.8269 -15.3258 -15.0467 -14.8236 -14.2665 -13.7094 -13.4304 -12.8733 -12.5942 -12.3152 -11.7581 -11.201 -10.6999 -10.1428 -9.9197 -9.6966 -9.1395 -8.5824 -8.3033 -8.0243 -7.4672 -6.9101 -6.353 -6.0189 -5.4618 -4.9607 -4.6817 -4.4586 -3.9575 -3.6785 -3.3994 -3.1203 -2.8412 -2.5621 -2.283 -2.0095 -1.4524 -1.1733 -0.8942 -0.6151 -0.336 -0.0569 0.2222 0.5012 0.7747" fill="rgb(0,0,0)"> During the combustion of gasoline, energy is ......1...... . </svg:tspan><svg:tspan font-family="g_font_9" font-size="1px" y="17.8798" x="-25.6771" fill="rgb(0,0,0)">●</svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="17.8798" x="-25.0703 -23.7363 -23.0132 -22.4561 -22.122 -21.8989 -21.3418 -20.7847 -20.5057 -20.2266 -19.6695 -19.1124 -18.8334 -18.2763 -18.0532 -17.4961 -16.995 -16.7159 -16.3818 -15.8247 -15.6016 -15.1005 -14.5994 -14.3763 -13.8752 -13.5962 -13.0391 -12.7656 -12.4866 -11.9855 -11.4284 -11.2053 -10.9262 -10.3691 -10.035 -9.8119 -9.3108 -9.0318 -8.4747 -7.9736 -7.7505 -7.1934 -6.9143 -6.6353 -6.0782 -5.5211 -4.964 -4.6299 -4.0728 -3.5717 -3.2927 -3.0696 -2.5685 -2.2895 -2.0104 -1.7313 -1.4522 -1.1731 -0.894 -0.6149 -0.0578 0.2213 0.5004 0.7795 1.0586 1.3377 1.6168 1.8958 2.1693" fill="rgb(0,0,0)"> During the electrolysis of sulfuric acid, energy is ......2...... . </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="19.0328" x="-31.4882" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="20.1858" x="-29.553 -28.6075 -28.05 -27.8265 -27.325 -26.7675 -26.4885 -25.765 -25.2075 -24.873 -24.3155 -23.814 -23.535 -23.0335 -22.476 -21.6415 -21.084 -20.8605 -20.303 -20.0235 -19.466 -19.1925 -18.635 -18.0775 -17.52 -17.0185 -16.7395 -16.182 -15.903 -15.3455 -14.788 -14.2305 -13.957 -13.3995 -12.842" fill="rgb(0,0,0)">Which words complete gaps 1 and 2? </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="21.3388" x="-31.4882" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="22.8634" x="-28.2574 -23.5012 -22.9437 -16.0008 -15.4433" fill="rgb(0,0,0)"> 1 2 </svg:tspan></svg:text></svg:g><svg:g transform=""><svg:path d="M 70.68 329.6 L 71.16 329.6 L 71.16 329.12 L 70.68 329.12 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 70.68 329.6 L 264.06 329.6 L 264.06 329.12 L 70.68 329.12 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 263.58 329.6 L 264.06 329.6 L 264.06 329.12 L 263.58 329.12 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 70.68 329.12 L 71.16 329.12 L 71.16 309.26 L 70.68 309.26 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 99.06 329.12 L 99.54 329.12 L 99.54 309.26 L 99.06 309.26 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 181.26 329.12 L 181.74 329.12 L 181.74 309.26 L 181.26 309.26 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 263.58 329.12 L 264.06 329.12 L 264.06 309.26 L 263.58 309.26 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:text transform="matrix(10.9755 0 0 10.98 81.12 291.9803) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_3" font-size="1px" y="0" x="0 0.7214" fill="rgb(0,0,0)">A </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="0" x="3.362 3.919 4.142 4.643 5.2 5.757 6.036 6.593 7.15 7.429 10.8623 11.4193 11.6423 12.1433 12.7003 13.2573 13.5363 14.0933 14.6503 14.9293" fill="rgb(0,0,0)">given out given out </svg:tspan></svg:text></svg:g><svg:g transform=""><svg:path d="M 70.68 309.26 L 264.06 309.26 L 264.06 308.78 L 70.68 308.78 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 70.68 308.78 L 71.16 308.78 L 71.16 287.78 L 70.68 287.78 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 99.06 308.78 L 99.54 308.78 L 99.54 287.78 L 99.06 287.78 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 181.26 308.78 L 181.74 308.78 L 181.74 287.78 L 181.26 287.78 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 263.58 308.78 L 264.06 308.78 L 264.06 287.78 L 263.58 287.78 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:text transform="matrix(10.9755 0 0 10.98 81.12 270.9803) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_3" font-size="1px" y="0" x="0 0.7214" fill="rgb(0,0,0)">B </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="0" x="3.362 3.9194 4.1428 4.6442 5.2016 5.759 6.038 6.5954 7.1528 7.4322 11.1443 11.4237 11.9811 12.4825 13.0399 13.5973 13.8763 14.0997 14.6517" fill="rgb(0,0,0)">given out taken in </svg:tspan></svg:text></svg:g><svg:g transform=""><svg:path d="M 70.68 287.78 L 71.16 287.78 L 71.16 266.78 L 70.68 266.78 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 99.06 287.78 L 99.54 287.78 L 99.54 266.78 L 99.06 266.78 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 181.26 287.78 L 181.74 287.78 L 181.74 266.78 L 181.26 266.78 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 263.58 287.78 L 264.06 287.78 L 264.06 266.78 L 263.58 266.78 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:text transform="matrix(10.9755 0 0 10.98 81.12 249.9803) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_3" font-size="1px" y="0" x="0 0.7214" fill="rgb(0,0,0)">C </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="0" x="3.6408 3.9202 4.4776 4.979 5.5364 6.0938 6.3728 6.5962 7.1482 10.8603 11.4177 11.6411 12.1425 12.6999 13.2573 13.5363 14.0937 14.6511 14.9305" fill="rgb(0,0,0)">taken in given out </svg:tspan></svg:text></svg:g><svg:g transform=""><svg:path d="M 70.68 266.78 L 71.16 266.78 L 71.16 245.78 L 70.68 245.78 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 99.06 266.78 L 99.54 266.78 L 99.54 245.78 L 99.06 245.78 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 181.26 266.78 L 181.74 266.78 L 181.74 245.78 L 181.26 245.78 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 263.58 266.78 L 264.06 266.78 L 264.06 245.78 L 263.58 245.78 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:text transform="matrix(10.9755 0 0 10.98 81.12 228.9803) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_3" font-size="1px" y="0" x="0 0.7214" fill="rgb(0,0,0)">D </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="0" x="3.6408 3.9205 4.4782 4.9799 5.5376 6.0953 6.3743 6.598 7.15 11.1409 11.4206 11.9783 12.48 13.0377 13.5954 13.8744 14.0981 14.6501" fill="rgb(0,0,0)">taken in taken in </svg:tspan></svg:text></svg:g><svg:g transform=""><svg:path d="M 70.68 245.78 L 71.16 245.78 L 71.16 224.24 L 70.68 224.24 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 70.68 224.72 L 99.06 224.72 L 99.06 224.24 L 70.68 224.24 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 99.06 245.78 L 99.54 245.78 L 99.54 224.24 L 99.06 224.24 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 99.54 224.72 L 181.26 224.72 L 181.26 224.24 L 99.54 224.24 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 181.26 245.78 L 181.74 245.78 L 181.74 224.24 L 181.26 224.24 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 181.74 224.72 L 263.58 224.72 L 263.58 224.24 L 181.74 224.24 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 263.58 245.78 L 264.06 245.78 L 264.06 224.24 L 263.58 224.24 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 263.58 224.72 L 264.06 224.72 L 264.06 224.24 L 263.58 224.24 Z" stroke-miterlimit="4" stroke-linecap="butt" stroke-linejoin="miter" stroke-width="0.75px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:text transform="matrix(10.9755 0 0 10.98 49.62 214.0403) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_2" font-size="1px" y="0" x="0" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="1.1475" x="0" fill="rgb(0,0,0)"> </svg:tspan></svg:text></svg:g></svg:g></svg:svg>
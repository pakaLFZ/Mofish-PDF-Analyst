<svg:svg xmlns:xlink="http://www.w3.org/1999/xlink" xmlns:svg="http://www.w3.org/2000/svg" version="1.1" width="595px" height="842px" viewBox="0 0 595 842"><svg:g transform="matrix(1 0 0 -1 0 842)"><svg:defs ><svg:style type="text/css">@font-face { font-family: &quot;g_font_3&quot;; src: url(data:font/opentype;base64,AAEAAAANAIAAAwBQT1MvMmLSWIkAAADcAAAATmNtYXAC9eNxAAABLAAAAHxjdnQg+z6j2gAAAagAAAdaZnBnbQjouigAAAkEAAAF12dseWaWaQK/AAAO3AAAQU5oZWFk5yaHjQAAUCwAAAA2aGhlYRJ+FiYAAFBkAAAAJGhtdHhZvsAMAABQiAAANXRsb2NhA1paJAAAhfwAADV4bWF4cBVHAbMAALt0AAAAIG5hbWXwxPICAAC7lAAAAmpwb3N0AAMAAAAAvgAAAAAgcHJlcPFK5RYAAL4gAAAR0gAABAABkAAFAAAEAAQAAAAEAAQABAAAAAQAAGYCEgAAAQEBAQEBAQEBAQAAAAAAAAAAAAAAAAAAAAA/Pz8/AEAAIAB5CAACAADMCCQEAgAAAAAAAQADAAEAAAAMAAQAcAAAABgAEAADAAgAIAA5AFAAVQBZAFsAaQBwAHcAeeAA//8AAAAgAC4AQQBSAFkAWwBhAGwAcgB54AD////j/+P/4//j/+P/4//j/+P/4//jIAMAAQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAW6ABwFugAcBacAHAQmABwAAP/kAAD/5AAA/+T+af/kBboAHP5p/+QC6gAAAR0AAAEdAAAAAAAAAAAAsgCsANcBKAEgALMB+gAXAPgBGQExAEkABAD3AAMArwD9AJUAFABUAJYBEgAkABYAVQBJAQQBGQErAIwBm/92/+kAPQCSAKL/twGC/6oAFgCPAMYA+AAcAN4EAQA3AE4AVQBVAGUA6QPlAFn/mgAIAIcACwA7AFIBFgBhANYA1gD1AAAAkwCUAL4BfP/4AAQAFACCAJIAPABBAEH/wf/8ACoAjASQBdgJtQCRALsBBv9j/2kAHgAiAIoCK//W/98AJgBZAKMArAEEASsBwARIACEAawCFAJgBGQPGAGsAlQCkAP4BDAJdA0MFvwAAAEkAVgBuAHcAigCqAMoBEgFQBdgF8P97/+cABgATACgAYQBpAOkBNQFNAqUEDP8+/9oAWwC5AMgBGQEZARkBwARbBKcFW/4//53/wgAVALcBCgG8AcEFMgWO/YH/of+uAAwAJgAxAD0ATgBWAGIAgwDBAMkA8QDyAn//fwBIAFMAdwDFAR0BIAEmASgB1gIZAn4CfgPTAC4AQQBdAGsAdQCfALAAsgC6ALsAvQDWANsA4ADlARQBGwFKAWIBkQHyAgwCZALPA5sDtAPUBAEEqQAWACMAJQAqAHQApQC2AMwAzQDPAQUBIAEwAVABagFvAZcBnQHgArAC7AL3BAgEgwT7BP0FJv7g/vv/Tv/1ABgAGgBMAHoAfwCRAKMAswC0AM4A1QDyAPMA9gEQATgBaAGhAbAB4AHsAgkCIgJPAnAClgKlAq0DTgORA8EENQRCBGsEzQTaBYYFiwdhB/78pv6T/q3+0f+3/9EAAwAOABgAJgBGAGkAgQCPAKUAvwDTANUA2QDdAOIBGQErATgBOwFaAV4BaAFzAYgBlAGtAcUB0QHqAfICAAIAAgACIgI7AkQCTwJvAnICfgKCApMClAKlAs8CzwLQAtoC3QLrAvUDBQMiAzYDcQOhA7ADuAPQA+YEEAQmBC4EMQRPBFoE/wUyBTIFRwVTBagFqwXCBfAGPAZkBnAG6AeCB4QIzP0q/d7+AP5o/rD+s/+qAAgAWQB6AJEAngCiAK8AtAC7AMoAzADOANkA4AD0ARQBGgEhAScBKwE5AUYBSwFNAVcBXAFlAYIBhwGSAZgBmwGiAa4BxQHFAdECBwIiAisCQQJTAmECZQKEAocCjQK0ArQCugLJAtYC2ALtAvUDFwMjAysDMQNJA1oDWwNuA3EDdAN+A4QDkQORA6oDzwPTA+cD6APtBAgEFwQeBHUEegSZBKcEtATRBUwFbQVtBaIFvwXABdEF/AX8BgIGGgYcBi8GagaoBuIHBgc2B1AHiQfUB/MIcAEcASoBGgEgAAAAAAAAAAAAAAAAAhkACwAeAqoCFAR/Ae0AAAAdAQQADwCRACsBiAFTARIB8wA/A/4BaAEOBH8B7QNuAxUCGQQTAAAAAAZABLAAAAJ0AbsANQHFAH8GAgMBAAAE4ACyAdwC4ATDAj0A1QFgARkEpwNuBcoCIQCrBCYAkAK8ArsBQgC0AjwCVgKcAwAB5QGoAOUAawB4AJQBawFzAKsB7QE6AX0BNwF/ANQCFgNTAYQAPP+iAgQBCQFJAfAAbgMVAIEEZABeAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAATkA3ADp/p4EDQR8ASsAuACWAFkArADfAakA+gEF/+wAFwADAFUAYQAEAIwAowCFACgBIABdANYAfwEmARkBBAFsBs8AtAEGAAAHNwY+BHoA8AD5AOkFugQmBEIAAP/n/mkEngTj/zf/LQEgAQUBIACoAHQAaABHAPIA5QDZAL0AqABoAEcAXABIAAoAKAAyAEEAUABaAGQAfQCHAJH/sP+c/4P/ef9vAMsBIAD6ASwB+gGgANUAuABcADwAyADIAI8A2QGLALMARwAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAP5kAMAA6gEYASUBMgOwA+0FdgWQBaoFtAW+Bc0GMQB4AIQAmwDMAOIA9AEKASABYwDRAOoA9wEIAUIAGQAsADQAQQA4AEgAWABsAlkDvQBDARoAcADTACgANwBCAFAAWgBkAHMAeACCAIwAnAClAL0AzgDwARABXAC+ANgBAgEXASwBYwDqAQgAQQBLAFUAXwBzAKYBCQGDAbMAQQBkAB4AKgDrAPoBDgE4AnQALABAAIIAlgC2AMAAzADcAOYA8AD/AQoBIAEsATsBRAFWAWMA9wBXAGQBEAE2AFABsQAA/7YAOQBOAEQDzADlACQBEABCASIBpADwAGAA4AAOAB0AOQXjAQIALP5O/zgCaQO9ARYA/wAOAKAAVAAbAD0BcQBBAA8AUAD9ABUBTwA1/lIALADTAQMEsAHSALYAwACZAmX/hwN3/mwAywCpAFwAQAR2B0QAAEBBVEA/Pj08Ozo5ODc1NDMyMTAvLi0sKyopKCcmJSQjIiEgHx4dHBsaGRgXFhUUExIREA8ODQwLCgkIBwYFBAMCAQAsRSNGYCCwJmCwBCYjSEgtLEUjRiNhILAmYbAEJiNISC0sRSNGYLAgYSCwRmCwBCYjSEgtLEUjRiNhsCBgILAmYbAgYbAEJiNISC0sRSNGYLBAYSCwZmCwBCYjSEgtLEUjRiNhsEBgILAmYbBAYbAEJiNISC0sARAgPAA8LSwgRSMgsM1EIyC4AVpRWCMgsI1EI1kgsO1RWCMgsE1EI1kgsJBRWCMgsA1EI1khIS0sICBFGGhEILABYCBFsEZ2aIpFYEQtLAGxCwpDI0NlCi0sALEKC0MjQwstLACwFyNwsQEXPgGwFyNwsQIXRTqxAgAIDS0sRbAaI0RFsBkjRC0sIEWwAyVFYWSwUFFYRUQbISFZLSywAUNjI2KwACNCsA8rLSwgRbAAQ2BELSwBsAZDsAdDZQotLCBpsEBhsACLILEswIqMuBAAYmArDGQjZGFcWLADYVktLEWwESuwFyNEsBd65BgtLEWwESuwFyNELSywEkNYh0WwESuwFyNEsBd65BsDikUYaSCwFyNEioqHILDAUViwESuwFyNEsBd65BshsBd65FlZGC0sLSywAiVGYIpGsEBhjEgtLEtTIFxYsAKFWViwAYVZLSwgsAMlRbAZI0RFsBojREVlI0UgsAMlYGogsAkjQiNoimpgYSCwGoqwAFJ5IbIaGkC5/+AAGkUgilRYIyGwPxsjWWFEHLEUAIpSebMZQCAZRSCKVFgjIbA/GyNZYUQtLLEQEUMjQwstLLEOD0MjQwstLLEMDUMjQwstLLEMDUMjQ2ULLSyxDg9DI0NlCy0ssRARQyNDZQstLEtSWEVEGyEhWS0sASCwAyUjSbBAYLAgYyCwAFJYI7ACJTgjsAIlZTgAimM4GyEhISEhWQEtLEuwZFFYRWmwCUNgihA6GyEhIVktLAGwBSUQIyCK9QCwAWAj7ewtLAGwBSUQIyCK9QCwAWEj7ewtLAGwBiUQ9QDt7C0sILABYAEQIDwAPC0sILABYQEQIDwAPC0ssCsrsCoqLSwAsAdDsAZDCy0sPrAqKi0sNS0sdrgCNiNwECC4AjZFILAAUFiwAWFZOi8YLSwhIQxkI2SLuEAAYi0sIbCAUVgMZCNki7ggAGIbsgBALytZsAJgLSwhsMBRWAxkI2SLuBVVYhuyAIAvK1mwAmAtLAxkI2SLuEAAYmAjIS0stAABAAAAFbAIJrAIJrAIJrAIJg8QFhNFaDqwARYtLLQAAQAAABWwCCawCCawCCawCCYPEBYTRWhlOrABFi0sS1MjS1FaWCBFimBEGyEhWS0sS1RYIEWKYEQbISFZLSxLUyNLUVpYOBshIVktLEtUWDgbISFZLSywE0NYAxsCWS0ssBNDWAIbA1ktLEtUsBJDXFpYOBshIVktLLASQ1xYDLAEJbAEJQYMZCNkYWSwA1FYsAQlsAQlASBGsBBgSCBGsBBgSFkKISEbISFZLSywEkNcWAywBCWwBCUGDGQjZGFkuAcIUViwBCWwBCUBIEa4//BgSCBGuP/wYEhZCiEhGyEhWS0sS1MjS1FaWLA6KxshIVktLEtTI0tRWliwOysbISFZLSxLUyNLUVqwEkNcWlg4GyEhWS0sDIoDS1SwBCYCS1RaiooKsBJDXFpYOBshIVktLEYjRmCKikYjIEaKYIphuP+AYiMgECOKuQKnAqeKcEVgILAAUFiwAWG4/7qLG7BGjFmwEGBoATotLLECAEKxIwGIUbFAAYhTWli5EAAAIIhUWLICAQJDYEJZsSQBiFFYuSAAAECIVFiyAgICQ2BCWbEkAYhUWLICIAJDYEIASwFLUliyAggCQ2BCWRu5QAAAgIhUWLICBAJDYEJZuUAAAIBjuAEAiFRYsgIIAkNgQlm5QAABAGO4AgCIVFiyAhACQ2BCWVlZWS0AAAIBAAAABQAFAAADAAcAQrQCAf4GB7gCP0ATAAUE/gMACgcE/gEAGQgGBf4CA7wBJgAJAbABGAAYKxD2PP08ThD0PE39PAA/PP08EPw8/TwxMCERIRElIREhAQAEAPwgA8D8QAUA+wAgBMAAAAEAkwAAAawBGQADACRAFQI4AAoCJg8AHwAgADAABAAZBGd2GCtOEPRdTf0AP03tMTAzESERkwEZARn+5wAAAf/9/+cCOwXTAAMAOEAdAAEBSQIDFAICAwIBAAMACgHrAhoFA+sAGQSTbBgrThD0Te1OEPZN7QA/PD88hwUuK30QxDEwBwEzAQMBa9P+kRkF7PoUAAACAFb/5wQOBcAADgAgAJNAS3gKiAqnAaoHqgmnDrcJyAkIVhFZFlkaVh9nEWgWaBpnHwg5AjkGNgk2DUkCSQZFCUYNpwnLAskGxAnEDdkC2wbUCdQNERAYIBgCGLj/wEAlEhY0GKYIDR8PLw8CD0ASFjQPpgAFHdhPBAEEGiIU2AsZIdPCGCtOEPRN7U4Q9nFN7QA/7StxP+0rcTEwAV0AXV0BMhcWERAHBiMiABEQNzYXIgYHBhEQFhYzMjY3NhEQJiYCMtV4j5B31db++pB31TNQFh00TzMzUBYdNE8FwJi0/l/+YLaWAUkBpgGetpbpQVRt/v7+/sFAQVRsAQIBAsFBAAEAogAAAyYFwAAJAFZACWsCewKLAgMCBLgBKbNfBQEFuAJetwgJBQEADAkAuwFYAAIAAQJdQA0FAAQfBCAEsAQEBBkKugGnAaAAGCtOEPRdPE32PP08AD88Pzz0Xe05MTAAXSEhEQYHNTYkNzMDJv7nmtFuAQIw5AQjkEX/JMmGAAABADMAAAQMBcAAHQE/QF+1GLYauRvKBMcY0BjQGdAaCEMbQxxDHVYZmwSVGKoEphwIBhogACgGNxpIBEMYQxlDGggkGCQZJBoDFiYEVgSIGJwbnBycHaocqh0IEgAdEB0gHTEddh2EHZAd1h0IHbj/wEAWFBU0HQIQDA8dEAAgAAIgADAAQAADALj/wLMSFjQAuAKhswIBDA+4AVZAIx8MLwwCDEASFjQMphMFCdgWFgFPAAEAGh8P2BB3Ahke08IYK04Q9E307U4Q9nE8PE0Q7QA//Stx5D88/StdcTwREjkBETMrXUNcWLkAHf/AshE5Hbj/wLIPOR24/8BADhA5BAgQOQUIETkECBE5KysrKysrWbEGAkNUWEALCRsZGwIbEwEEEwAAERI5ERI5XVkxMAFdS1FYvQAb/+AAHP/gAB3/4Dg4OFkBcV1dXQERITYSNzY3NjU0JiMiBgclNiQzMhYVFAYHBgQGBwQM/CcQoOy+KzplWVhoCP7oGQEIxtn4R00z/vZHFgEF/vuUAQnbsT9XVV5lansc6MrqrmOzYkH0UCYAAAEATf/nBBsFwAApANlAMocVyRUCexyLHAKmA6kFpxS2A7oFthTaGN0ZCBYUAY0WjRcCIQoNAAQBFxMWIR8NEAwKuAEkQAxPDQFADY8NAg0NARa4AQJADx8TLxMCE0ASFjQTphsFAbgBVrUQBCAEAgS4/8BAMhIWNASmJw2wDMAMAgwMFhDYfx+PH58frx+/HwUf4AfYTyQBJBorFtgXdwHYABkq08IYK04Q9E3t9O1OEPZxTe30Xe0ROS9dAD/9K3HkP/0rceQROS9dce0BERI5ETkAERI5ERI5ERI5XTEwAXFdXQBdEyUWFjMyNjU0JiMiBzcWNjU0JiMiBgclPgIzMhcWFRQHFhYVFAAjIiRNARANclFXd3JSNksfcnhYSUhmC/79G23Dec99Z9N+l/7m0sf++gGFIWhuhHBqfBXlA2lXSlhkYCyFn1uEbIjBcxu8hcH+8OUAAgAmAAAERAXAAAoADQDfQDkMIA05CQwZDCsMUwxrDOIMBu0NAQYEFgQlBCgNSA1bDacNtw3GDQkBAggADAYNBwUKCw0HAAwMDQ24Aa5AGgMEFAMDBAMCDAQNAw0CBAoAB0ANwA3QDQMNuwEoAAgAAgG0tgAEBAAMDAC4AVi0BY8KAQq4AQJAEhAHnwe/BwMHGg8/An8CAgIZDroBTAFIABgrThDkcRD2XU30XTz9PAA/PxD0PP1dPAEREjkSOTkAERI5EjmHBS4rBH0QxA8PD7EGAkNUWEALLQw9DE0MzQzdDAUAXVkxMAFdXQBdKyERITUBMxEzFSMRAREBAn79qAJ87La2/vD+rwEn9gOj/F73/tkCHgH1/gsAAQBb/+cENQWmAB0BEEApCA4gDDcSRRJJGZkNng6XEtoOCRIRExIhESMShRIFAAQBDQoMDA0SERG4AqBAFg4NFA4ODRIKFCABMAFAAQNQAZABAgG4AVa1EAQgBAIEuP/AtxIWNASmGw0MuAJaQA0fCi8KAgpAEhY0CqYUuP/AQAsUFjQgFDAUQBQDFLgBq0AUEREfEC8QAi8QPxBPEAMQQBIWNBC4AqBAEw8PDgQPEOAH2NAXAUAXARcaHw64ASFAEg13AbzQAAFAAJ8ArwADABke07kBRwAYK04Q9F1xTe305E4Q9l1xTe30PAA/PBD9K11xPBD2XSv9K3HkP/0rceRdcRESOYcFLisOfRDEARE5ABESORESOTEwAXFdEyUWFjMyNjU0JiMiBycTIREhBzYzMgAVFAcGIyIkWwEYDHZNWHp5YXlg5JAC5/3uLF5iuwEEaY/+y/8AAXkdX2+PkIeHayEC+/75+S/+8Nm1jsLaAAIAV//nBCoFwAAXACMAvUA7agt1CIcIlxmnBacIqQ6qE7kOthG9E8ARzxMNFQU2EUQQeha1AtIQ0BQHuwDPAAIABAEHGBIQGyAbAhu4/8BAHhIWNBumDw0fIS8hAiFAEhY0IaY/CQFACdAJ/wkDCbgBT7OvAQEBuAEhQCIfBC8EAgRAEhY0BKYVBQHYAHce2E8MAQwaJRjYEhkk08IYK04Q9E3tThD2cU3t9O0AP/0rcfRd9l1x7StxP+0rcQEREjkAERI5XTEwAV0AXQEFJiYjIgYHNjMyEhUUACMiABEQADMyFgEUFjMyNjU0JiMiBgQP/vAKVENZexBpnLD7/vjP3v7iASrup9v9oX5RTmhwVFFwBFMeVFCg/Xz+9NTh/vABWQGJAZMBZLv86YmVeouPhX8AAQBXAAAEGAWmAAsAhrkABP/gQDEPETQKCxoLOgQ4CkgFVguqC74LzQvZCwohCwELAwcAHwsvCwIvCz8LTwsDC0ASFjQLugKgAAMBrLcCAgEEBwgMCLgBWLMvBwEHuAJgQA4CTwMBAxoNAQAZDNPCGCtOEPQ8EPZxPE30Xf0APzw/PBDt/StdcTwBERI5XTEwAV0rExEhFQYCAhchEhI3VwPBd/aBAf7xB+3GBKEBBcx1/kr+E8IBMAJ4+QADAFP/5gQXBcAAGAAkADABDbUwCB0fNCa4//hAbB0fNMcRxxPXBdcHBHUQdhSEEAMmACoMNgA7DEYATAxuBGMIZxFoFXcnhyeXDZgYpA2pGKkaph6nJ6YsqTC5GrceF3cThhOGFIcnBJcMAQyXAAEAHC6YDAEMKwmXAAEAJQMuQBIWND8uTy4CLroCjgAc/8BAEBYYNHAcgBwCoBwBHBwGEii4/8BACRIWNDAoQCgCKLgCjkANEg0/Ik8iAiJAEhY0IrgCjkAaBgUf2Al3K9hPDwEPGjIZ2AN3JdgWGTHTwhgrThD0Te307U4Q9nFN7fTtAD/tK10//V0rEBE5L11xK+1dKwEREjldERI5XQAREjldOV0xMAFxXQBxXSsrASYmNTQ2MzIWFRQGBxYWFRQEIyInJjU0NhMUFjMyNjU0JiMiBgMUFjMyNjU0JiMiBgFIbWPl09HnamB6f/7918iFnXa5X09QYF9OUWAad1lXcnRZZ2UDFy6hYKTW1qRmnyoxvHvL/ml82HfHAVFUXl9UT19g/T10gn12Z32OAAACAEH/5gQUBcAAFwAjANBAWDsRSxFlC3oIiQipBakIpg6mE7UAuQO1DrgRtBPFAMoRwBMRNBNWC1kNXxFSE2ATBhkFdxaZF90Q3xQFaBMBAAQBBxgSHxsvGwIbQBIWNBumDwUQISAhAiG4/8BAEBIWNCGmMAkBTwnfCfAJAwm4AU+zoAEBAbgBIbUQBCAEAgS4/8BAGxIWNASmFQ0Y2E8SARIaJQHYAHce2AwZJNPCGCtOEPRN7fTtThD2cU3tAD/9K3H0XfZdce0rcT/tK3EBERI5ABESOTEwAXFdAHFdEyUWFjMyNjcGIyICNTQAMzIAERAAIyImATQmIyIGFRQWMzI2XQEQClRFV3oRap+t+wEJzd8BHv7W76zUAl59Uk5ncFRRbwFTHlNQoPx7AQvW3wER/qf+df5u/py3AxyIlnuMjoWAAAIAAAAABb8FugAHAAoBQbkAB//YQAk3OTQGKDc5NAe4/8BACSg1NAZAKDU0B7j/2EBQISc0BighJzQpACoEKgUoCi8MOAA3BT8MagBqAmUDZgVoCGcK6AMPSgYBAggJAQMKCQkEBwkBASAABxQAAAcGCQQEIAUGFAUFBggKQBodPgq4/8BACxodNAolAgMDBgQJuAG8QA4GBwIFBAQBAAgMFxcaALgCYUALHwEBIAEwAYABAwG4AiRACR8JATAJgAkCCboCJAAEAmFACSAFAQUZC15jGCtOEPRdTf0Z9l1x9F1xGP1ORWVE5gA/PDwQPD88Te0REjkvPP0rKzyHBS4rh33Ehy4YK4d9xAcQPDyHxMSxBgJDVFi0CTQJDTQAK1kxMAFLsAtTS7AeUVpYuQAD//6yCAQKuv/+AAf//LEGBDg4ODg4WQFxXSsrKysrKyEhAyEDIQEhEwMDBb/+voD9tnn+xgI7ATkqysYBTf6zBbr8igIg/eAAAAMAlgAABWIFugATACAALADYQD93KgFoDngq5gT2BAQJIRUJBigsISUWEh8VTxUCMBWvFQIVFRQjIiUSEwggFCUBAAIbJ3AGgAYCBksoJ68MAQy4/8CzCQs0DLgCjEAhMC5ALlAuYC5wLoAukC6gLgggLjAuAi4UIiAAIBMwEwITuAKLsy0xUxgrThD0XTxN/TxNEF1x9itxTe30Xe0APzz9PD88/TwROS9dcUNcWLkAFf+Ash05Fbj/wLIaORW4/4CxEzkrKytZPP08ARESOQAREjkxMAFLsAtTS7APUVpYsQogOFkBXQBdEyEyHgIVFAYHFhYVFAYGBwYFIQERMzI3NjY1NCYnJiMDESEyNzY2NTQmJiOWAkquq4dab1+GkF2hdkr+5f4NASjCrSpMV0tKLNGqARKgK0JTQHnKBbodXJlfZ6wrJ7x/ZL1xDQgCBMb+rQUJV0dEVQkF/bn+eAkMXU5CXCoAAAEAYf/nBV4F0wAaANZAToYJiRSJFp8AmAbHCdQD1Av1AwklCSgMKA0pFCkWdQV1CYYFCAcTBxcXExcXKQIqAyUFBygFmQWXCckDxQsFPwFPAQIBUhAAAeAA8AACALj/wLMRGDQAuP/AswoNNAC4AVpAFxgtBAgOQA4SNA5LXw8BTw8BD0AVGDQPuAEoQCISLQoDD+8OVgDvAAFPAQIBGjAcARwVJ6AHAQ8HHwcwBwMHuAKMsxt+UxgrThD0XXFN7U4QXfZdTe307QA//fQrXXHkKz/99CsrXXHkXTEwAF0BXV1dAQUGBCMgABEQACEgFxYXBSYmIyIGERAWMzI2BD8BH0L+zez+3P6IAXoBNAENqGQy/tsapXajy8igdqoCG1vw6QGPAVoBbgGVn16wRnKE6v76/urslgAAAgCUAAAFYQW6ABAAHwB/QDMoBSgKRxdlBGUMBSoXORdIFlkWaBYFORc2G4cbmQWWCwUfESUBAAITEiUPEAgZJ68HAQe4/8CzCQs0B7gCjEATgCEBICEwIQIhERIgACAQMBACELgCi7MgMVMYK04Q9F08Tf08TRBdcfYrcU3tAD88/Tw/PP08MTAAXXEBXRMhMhcWFhIVFAcGBwYHBiMhAREzMjc+AjU0JiYnJiOUAh23YIG4YC03Zk2DYqT90wEo3Xw3SF88PGxTPrUFuhwmwv7nzrWDoGNLKh8Ewvw1DhJWxaqqtmYSDgAAAQCVAAAE8AW6AAsAkEA9CAUEBwglBhIfBQEwBa8FAgUFCQMEJQIBAgoJJQsACAcGSwMCSAoACwELGiANMA1ADQMNBAkgASAAMAACALgCi7MMMVMYK04Q9F08Tf08ThBd9l08TfQ89DwAPzz9PD88/TwROS9dcUNcWLkABf/Ash05Bbj/gLIaOQW4/4CxEzkrKytZPP08AwUQPDwxMDMRIRUhESEVIREhFZUEP/zpAuD9IAMzBbr4/rv3/nH3AAEAlwAABIQFugAJAHJAPwgFBAYFJQcgCDAIvwjfCAQvCJAIAggIAAMEJQIBAgkACAc/Bk8GAgZSAwACAQIaIAswCwILBAkgASAAMAACALgCi7MKMVMYK04Q9F08Tf08ThBd9l08TfRdPAA/PD88/TwSOS9dcTz9PAMFEDw8MTAzESEVIREhFSERlwPt/TsCZP2cBbr4/qX4/ZEAAAEAYv/nBb0F0wAgANhARjgeSx5WB3YIdgyFCIQMhReEGwkGFwYbEhcSGygRKBgoGigeCEgLWwRUCVoLagR7BHoYdBq2DrYQxw3GENcQ5xAOAxwGIAC4/8BAHxo5HwABACUCAQEWHC0GCRJADhI0EktPEwETQBUYNBO4AShAKhYtDwMAAQEgGV8TARMnElYCHyAgAwIaICIwIgIiGSegCgEPCh8KMAoDCrgCjLMhfp8YK04Q9F1xTe1OEF32PE39PBD07XEREjkvPAA//fQrXeQrP+0ROS88/XErPBESOTEwAF0BXV0BNSERBgQjIiQCNTQSNzYzIAQXBSYmIyIGFRASMzI2NzUDPwJ+Xf6fteb+qqzAuY3SAREBMyz+2h+rgMLl6Lxdu0MCG/f9uFqJwQFn0+UBZF9J5co3bH328v77/vtJNLoAAQCWAAAFKgW6AAsAo0AlCQQFCgMCCQolBBKvAwEDAwAGBQUCAQIHCAgLAAgFCCAGzwcBB7gCi0AiQA1QDWANA3ANgA0CIA0wDaANwA0EDQILIAEgADAAwAADALgCi7MMMXUYK04Q9F08Tf08TRBdcXL2XTxN/TwAPzw8EDw/PDwQPBI5L11DXFi5AAP/wLIdOQO4/8CyGjkDuP/AsRM5KysrWTz9PAMFEDw8EDw8MTAzESERIREhESERIRGWASgCRAEo/tj9vAW6/b8CQfpGAoH9fwABAIwAAAG0BboAAwBvuQAF/8CzMjQ0Bbj/wLMjJTQFuP/AQD8UFzQABUAFUAWABeAFBR8FYAVwBfAFBIAFAQIBAgMACAID2QEAALAA4AADwADwAAIgADAA0ADgAAQAbgQxnxgrThD0XXFyPE39PAA/PD88MTABXXFyKysrMxEhEYwBKAW6+kYAAQAj/+cDzQW6ABIAWkAkaQinDQJUCWYJaQ1pEGkRehCJEAcKSAuBDy0HCQEAAgASIAECuAKLQBJwFAEwFAEUC+8fCgEKGRP9dRgrThD0XU3tTRBxcfY8Tf08AD88P/305DEwAF0BXQEhERQHBgYjIiYnJRYXFjMyNjUCpgEnICviudnqAQEXBSAwYmNSBbr8YLZigJvz6yB+NE9xsgABAJkAAAXDBboACwGRQBoIBgESEgoKBQMCAwQGBgcJCgkICgUJCAkKCLgBt0ArBwYUBwcGAwQEIAUKFAUFCgoJAwMGCgMJAwgLBgYHBQQEAgECAAsLCAcIBLgCZLIFSAi4AmRAEgcaIA0wDQINAgsgASAAMAACALgCi7MMMWMYK04Q9F08Tf08GU4QXfYYTe307QA/PDwQPD88PBA8GRI5LwEREhc5ABIXOYcFLhgrBH0QxIcFLhgrCH0QxIcIEDwIxAMIEDwIPLEGAkNUWLUJIAsNNAO4/8qyCCc0ACsrWTEwAENYQBkmBicJkASYBqAEsATABAeEBqgE6AT2BQQJuP/gszdSNAm4/8BAJDdSNCUGPQp0A4YDmQOZCZoKqgO6A8kDCsED0AP8CgM9CkIDAnJxXSsBK3FdWUNcWLkABv/osxILPwa4/+hAEw8LPwQwDRY/BDAMFD8EIAsSPwO4/9CzDxk/A7j/0LMOFz8DuP/Qsw0WPwO4/9CzDBQ/A7j/0LMLEj8DuP/Qsg4TPwArKysrKysBKysrKytZAV0zESERASEBASEBBxGZASgCVgGO/dgCRv6B/m3wBbr9dQKL/cX8gQKw9f5FAAEAnQAABKUFrgAFAD1AGlAHAQIBAgQDJQUACAQFGgcCAyABIAAwAAIAuAKLswYxuRgrThD0XTxN/TxOEP48AD88Tf08PzwxMAFdMxEhESEVnQEoAuAFrvtJ9wAAAQCRAAAGGQW6AAwCGEALCwMmCCYLAwQDAQO4/4BACRw6NAogOjs0Cbj/4LM6OzQJuP/gQKQcLjQKIBwuNAYJCArjCewKBAQJCgoTAhwEEAkfCiMCLAQgCS8KZwJoBGUJagp3AngEpAmqCrUJugr2CfoKFp8EkAmfCsYJyQrXAtgE1gnZCucC6ATlCeoKDXcJeAqDAowEgwmMCpACB1gLZQJqBGcJaAp2AnkEB0QCSwRECUsKVwhXCVgKBxgKLw40AjoENAk7Cj8OBwMCDAQGCQkKFQIaBBcJB7EGAkNUWEAfAgQDCgkFDAcHMgYODDIAAAMQAwIIUAgNNAtQCA00A7j/gEAOCw00CEAOJzQLQA4nNAO4/5xAEA4nNAMLCAMBAAQBAgcKAAgAPzw8PzwREhc5KysrKysrXQEv7RDU7RESFzkbuP87QC0DCgkgBAgJCTIDBBQDAwQCCwoKMgMCFAMDAgsIAwMMBAICDAoKCQkHCB8OAQ64AQ2zBwYFBLoCOAAF/8CzW100Bbj/wEAXU1Q0BTIHQAd/CAEIvX8DAQO9CyALDAK4AjhAEgEAAEBbXTQAQFNUNAAyHwwBDLgBDbMNMXUYKxD0ce0rKxA87hA8GhkQ/XH9cTwaGBD9KyvuEDwQ5HEAPzwQPBA8PzwSFzmHBS4rh33Ehy4YK4d9xCtZMTABS7ATU1i5AAj/4LELIDg4WQFdXV1dXV1xcisrKysAK3FdMxEhAQEhESERASEBEZEBuwEKAQcBvP7t/t3+4/7eBbr8GAPo+kYEgvt+BIL7fgABAJgAAAUjBboACQHOQA4JAwYIGQMXCAQSCAIDA7j/ALMSCz8DuP/As1tdNAO4/8BAKlNUNAMyBwgUBwcIAwgCAgcDCQQCAgkHCAMEQFtdNARAU1Q0BDIGzwUBBbgCi0AZQAtQC2ALA3ALgAsCoAvACwIgCzALAgsICbj/wLNbXTQJuP/AQA5TUzQJMgEgADAAwAADALgCi7MKMXUYK04Q9F08Tf0rKzxNEF1dcXL2XTxN/SsrPAA/PD88ARESOTkAEjk5hy4rKysrh33EsQYCQ1RYuQAD/+BACQ4nNAggDic0A7j/wLcJDTQIQAkNNAArKysrWTEwQ1i5AAP/gLYLNQiACzUDuP/AQD0aLjQIUxouNAUDFgMyA0ADBEYDhQiQCKAIsgjkAwbEA88I2ggDIAMvCDQDOwhPCJIDnwigA68IsAO/CAsHuP/AQAkzNTQCQDM1NAe4/+BADS8yNAIgLzI0AgcUNQe4/5dACSEuNAJUIS40B7j/wEBGHiA0AlQeIDQIAgcHGAIDFwcsAicHOwIzB04CQAdcAlYHCRQCGwdNAkUHmgerB8sC2QLoAucH+QILJwIoB0oHeAeIB6wCBgFdcXJyKysrKysrKysrAF1dcXIrKysrWQBdMxEhAREhESEBEZgBIAJYARP+1/2xBbr8LQPT+kYDvPxEAAACAFn/5wXnBdMADwAbAKJAVZcFlwiYDJgOBAgBBw4IDwcYJxh4CXcSB3cReBWGBIkIiQyGDoUSiRSIFYgXiBiGGgwHEggUBxoVEhoUGhgVGgcTLQ0JGS0HAxYnrwoBAAoQCiAKAwq4AoxAIDAdQB1gHXAdgB2gHQYgHfAdAh0QJ6AAAQ8AHwAwAAMAuAKMsxx+wxgrThD0XXFN7U0QXXH2XXFN7QA/7T/tMTABXV1xAF0TNDc2Njc2MyAAERAAISAAARQSMzI2NTQmIyIGWUMyrWeJswFEAYX+fv69/rn+fgEx5rGx4923t+AC1OCYcLIrOv5u/pr+nf5vAY8BaPn+/////Pj7AAACAJUAAAT4BboADwAbAHdAJQYFuRS5GANHBQFnBdYFAhIRJQ0ODgAbECUCAQIPAAgWJ68HAQe4/8CzCQs0B7gCjEAWHx0wHWAdcB2AHQUdEA8gASAAMAACALgCi7McMVMYK04Q9F08Tf08TRBx9itxTe0APzw/PP08EjkvPP08MTAAXXEBXTMRISAXFhYVFAYGBwYjIxkCMzI2NjU0JicmI5UB2wEOUn6qYpdOasnBoq92Q15INaAFuhYh3a+HuGkRFf3XBML+YC5iQVBoDQoAAgCWAAAFvAW6ABUAIQD4QII5D0kPVwdqC2oMqgmnDqAjtg7YCQoGCAYKFwgWCjYORg5GDwcIEAkRFA4UDxQQNg42D0cPdQ55ENMKC3gJeBl2HYgJiBmGHQYJFhQJDA8OUw51DoQOlA6jDgUOIA0MFA0NDA8MFQ0XFiUTEBQBYBSgFAIUFAAgISUCAQINDg4VAAgOuAG8QCcADRANAg3UGyegBrAGwAbQBgQGh3AjASAjMCMCIyEVIAEgADAAAgC4AouzIjFjGCtOEPRdPE39PBBdcfZd7fRd7QA/PDwQPD88/TwSOS9dcTz9PAEREjk5hy4rXQ59EMQBETkAERI5MTAAXQFxXV0zESEyFhYVFAYHFhYXEyEDLgIjIxERMzI2NjU0JicmIyOWAm/r1YDCwWB9arP+ntZyVF5mPNvVajxPSCS05wW6T8qCpdccOIar/uIBP6tZIf2cA04kWEJKWwwFAAABAEr/5gTyBdMALAHQQD25EbgdtijGLAQHEwcVFxMXFRgrZQVlKHQGeA10KNkM1iMMWQpVDlUiWSNoDGYSZyFpKGcsdx2GHZYhDBIjuP/gsx4fNCO4/+BAZRkaNFEiUSPBIsEjBHEicSOBIoEj4SLhIwYrCioNJCIkIzkNNCNLCksNRCJDI2oNZSN5DXoiiQ2KIqYKpw2oIhMJCgkNBiIGIxkKGQ0WIgciIwoNBAEXVhhAGSA0bxgBbxifGAIYugJlABv/wEAMGjkfGwEbLRQDAEgBuP/AQEkaIDQwAUABUAFgAZABoAGwAcABCAHuBEAaORAEAQQtKgkY7/8XARdAExc0F0sHJyYaLh8noBCwEAIQSwHvESAAMAACABkt0lMYK04Q9F1LU1ixAEA4WU3t9F3tThD2Te30K3LtAD/9cSv0XSvkP/1xK/RdcivkEhc5XV1xcisrQ1xYuQAi/+CzGx0+I7j/0LMbHT4juP/jshM5Irj/4LITOSO4/8myEjkiuP/QQA8SOQ0gEjkKIBI5CiAPOSK4/+hADgw5DSANOQoYDTkKGBM5KysrKysrKysrKysrK1mxBgJDVFhAFToKOg01IjUjSwpJDUMiRiOmCqkiCgBdWTEwAF1xAV0TJRYWMzI2NTQmJyYnJicmNTQ2NjMgBBcFJiYjIgcGFRQXFgQWFhUUBgQjIABKASAan4ePkT1MNLnuYId/76kBFAEXB/7YE319gUkvLDgBsM91jP8Av/7q/tYB3RyRiHlRNEkbEi47VnmucMNm8soNcWM1Ijk0JS9mbb2LftxrAQEAAAEALAAABLkFugAHAHJAIy8JMAQwBVAJcAmACZAJBwYBBQIlBAMCBwAICRcXGgR/BQEFuAEtQAoGByABMAB/AAIAuAEtQBEDDlACcAKAApACBAIZCP2sGCtOEPRdS1FYsQJAOFk8TfRdPP089F08RWVE5AA/PD88/Tw8PDEwAV0hESE1IRUhEQHf/k0Ejf5OBML4+Ps+AAEAk//nBSQFugAZAIpAOAcIBwkHEBcIFglHCEcJB1cJVhCWEJcRmBWbFqcQtxbXFeUG9gYLDQwMAQACByUTCQwLIA3PDgEOuAKLQCJAG1AbYBsDcBuAGwIgGzAboBvAGwQbAQIgACAZMBnAGQMZuAKLsxoxdRgrThD0XTxN/TxNEF1xcvZdPE39PAA/7T88PBA8MTABXXETIREUFxYWMzI2NjURIREQDgIjIiYmJyY1kwEoCxOPfH6AGgEoMIHYrtLZfhQdBbr85r04Wm1nlq4DK/z+/vjalllhm1V+9gAAAf/9AAAFWAW6AAgAxbkABP++QD4LNcAKAQQDBAUDBwQFBAMFAQQDBAUDIAIBFAICAQQFBAMFIAYHFAYGBwEEBwMGCAcEAQMCAwkEAAUKCAFWB7gCZ0ALBgYFBQMDAgIACAq7AhcACAAGAhe1BwcIIAACuAIXtwEBIAAwAAIAuAJmswleYxgrEPZdPBkQ5BgQ/TwZEOQYEOQAPz88EDwQPBD25AEREjkSORE5ABEXORESFzmHBS4rCH0QxIcFLhgrCH0QxAcIEDyHCBDEMTABXQArIREBIQEBIQERAhb95wFbAVkBUgFV/eUCaQNR/bwCRPyt/ZkAAQCS/mMChAW6AAcAUEAyBjAFQAUCBTcAAz8ETwQCBDcBEAASAwIGAgcEBRAHAQf0BZsAACABMAHQAQMBYAhnfBgrEPZdPBDt7V0QPBA8PBA8AD8//V08EP1dPDEwExEhFSMRMxWSAfLn5/5jB1fd+mPdAAACAEn/6AQuBD4AIwAyAXFAaAcaCBwFHRYaShtIHEkl2xDfEQk2GUYZVyZmGWcmhiaSGZMaphq5G8cayBsMBgYNFRYGGRYnBikVWRl3AoYCpga1BsYGDL802RACHSQyMREsDSRAKy40JEAiKDQkQBkdNG8k/CQCJEYduP/AQDAODzQ9HQEAHRAdsB35HQQdHSwBMwBADg80DwAfAAIAVSFAHBE/IUAbED8hQBgaNCG4AnS1BAcMDQosuP/AsxwRPyy4/8CzGxA/LLj/wLMYGjQsuAJ0QEAUCx4xJggpCSgNWR8MnwwCHwwB/wwBDEAOFjQMGk80ATRgAAEAjjABAQEzKSFfFwHfFwFPF18XbxcDFxkzaUEYK04Q9F1xck3t9HHtXU4QXfYrXXFyTe305P08AD/tKysrPzw//SsrK/RdK+QSOS9dcSuxBgJDVFiyLx0BcVntsQYCQ1RYuQAk/8C3Gx00VCRkJAJdK1ldKysrERI5Aw4QPDw8MTABcV0AXXEBJzY2MzIWFhUDFBYXISYnJicGBiMiJjU0NjY3Njc1NCYjIgYBBgYHBhUUFjMyNzY3NjUBZf8r0s+8uEsDGyX+6gsQBwNIpF2kvVabksVMUG9LVAFeNuokN1hETEUzEAsC4i6alFmJt/64jIVMHDcZCEZGsohajUscJSAcUUU7/tISMhgnPDtWMiY3JGUAAgCH/+gElAW6AA8AHACduQAS//hAMQs5NxtHGwISVgZWClYWVhhZHPcHBjUEOw07EzUbRQRLDUsTRRuUB5kJCgwOAQIBABq4AnSyBQcUuAJ0QBMLCw8AChchCBpwHgEeECkCAyYPuAEpQAwBcACAAAIAGR0/QRgrThD0cTxN7f085k4QcfZN7QA/PD/tP+0/PDEwAHFdAV1DWEALZgZmCmYWZhhpHAVdWQBdKzMRIRE2MzISERAAIyImJxUTFBcWMzI2NTQmIyIGhwEZgrLC/v79uVuxQBI0SXldg4RnZYYFuv3wlP7n/vn+8P7aW1mcAiqlT3Cfq7ahnQAAAQBV/+gEPwQ+ABkA4UBRWA9ZElkWaA9pEmkWfRh5GZcClwzGEMYY1xDWGOkG6QjpE+kV+AYTOBM4FUoSShZGGFkMaQwHOhI3FjcYA3cFdw+HBYYPiRmoEqcWuRK2FgkOuP/AsxgbNA64/8C1EhQ0DjMNuP/AsxkeNA24/8CzDxE0DboBBAAKAnRAEhELAEAYGzQAQBIUNAAzkAEBAboBAQAEAnRAIBcHAUASFDQBIQAvDUASFDQNIU8OAQ4aGwchFBkaWEEYK04Q9E3tThD2XU3tK/TtKwA//fRd5CsrP/30KyvkKysxMABdcQFxXQEFJiYjIgYVFBYzMjY3BQYGIyIAERAAMzIWBDH+6w5jT2l9f2tQZhUBFCv0zen+6wEW7cLlAuwyU1SRqr2cW28vvsIBJgEEAQcBJacAAAIAVP/oBGEFugAPABwAkEAtElkGWQpZElYWVhhZHJgHmQn4CQlwHoAeAjoDNAw6FTQZSgNEDEoVRBmZCQkUuAJ0sgULGrgCdEAOCwcODwABAAoXKQ4NJgG4ASlADw8AGo8eAR4QIQgZHVg8GCtOEPRN7U4QcfY8Te39POYAPzw/PD/tP+0xMABdAXFdQ1hADWkGaQppEmYWZhhpHAZdWSEhNQYGIyIAERASMzIXESEBFBcWMzI2NTQmIyIGBGH++0GxWrf++/7CsoIBGf0SL0R6YYiEZ2SHnFtZAScBCAEOARmUAhD8cKpMbqWkt6GfAAIAQf/oBCcEPgAUABwBo7kAEP/4QEYLOZkJmg2WEKgFpwq7CbsNuBoICBQBSAJHBkYKTx6oDbYGthrHCsgM1grYDPgH9w0NHA8cFUAbHTQVQA4RNA8VvxXPFQMVuP/Asw8ePxW4/8CzDhc/FbgCjUAMDw4SUA5gDgIOGBIBuP/AthkbNAEzEgC4/8CzHSA0ALj/wLMiKTQAuP/AsystNAC4/8CzGBw0ALj/wEAPDg80oAABAAAQAAIAXxISuAJ0swQLEhi4AnRAJAsHACEBLxUhTw4BDhovHl8ebx6fHgQeDyEIQA0PNAgZHWlBGCtOEPQrTe1OEF32XU3t9O0AP+1DXFhAFBhAKBQ/GEAeDz8YQBsQPxhAHBE/KysrK1k//UNcWLkAEv/AsygUPxK4/8CzHg8/Erj/wLMbED8SuP/AshwRPysrKytZ9F1xKysrKytDXFi5AAD/wLISOQC4/8CyFzkAuP+wswkKPgC4/8CyQSE/KwArKytZ5CsREjldQ1xYQBQOQA8ePw5AHBE/DkAbED8OQA4XPwArKysrWS88/SsrcisrPAERMzEwAV1xAF0rAQUGBiMgJyY1EAAzMgADIRYWMzI2EyYmIyIHBhcC+gEYNumv/uuFaQEU0+0BEgb9QAOCYUJaJwN4Vlw8PAEBUi+aobWR3QEIASv+x/69fYtIAWx6f0NDcwAAAQAYAAAC5gXTABYAuEAyNgQBKgQgECARWQSAGAUIBL8YAhUWEQIUEhYRDhMPABAOEwEAEAIUCQgPCwFfC/8LAgu4AnRACgYBEQ8WAf8WARa4AnRAHhAAAAHwAAEABhMUCgkzPwhPCFAIAwgoEC8RXxECEbgBBEANDhMmAhRfAKAWwBYCFrj/wLYJDDQWGRd4uQJpABgrThD0K3E8Tfw8/Tz8XTz0XRnkABg/PD9dcTz9XXE8P/1dcTkyDw8PDzEwAXFdAF0TMzU0NjYzMhcHJiMiBhUVMxUjESERIxicOZl1eHMmQz49NdLS/uecBCZQhoRTJMQQOVFL3fy3A0kAAAIAVP5RBGAEPgAjAC8BTkBidx2HHQISDA1wMYYNgDEEIAEjAiMDMAEzAjMDQAFDAkMDWw9ZFFklVilWK1kvaw/4EfgTEjsNMxY7KDMsSw1EFksoRCzwDP0XCo4MAQwLDA0LKgwNJw4WFxUtDQwXFgQYJAG4/8C1GRs0ATMAuP/Asw4RPgC4/8CzCww+ALj/wLMoKjQAuP/AsyMlNAC4/8CzMTQ0ALj/wEAJFRs0YAABAF8FuAJ0sh8PJ7gCdLIOCi24AnRACxUHGBkGKikLJhoYuAEpQAkZGRoajzEBMQG4AbhACgAzJCESGTBYPBgrThD0Te307U4QcfY8TRDtEP3kAD88P+0/7T/99HIrKysrKyuxBgJDVFi5AAD/wLMOETQAuP/AsgkMNCsrWeQrARESFzkAERI5ORESOTkHCBA8MTAAcV0BXXFDWEANaQ9pFGklZylmK2kvBl1ZAF0XBRYXFjMyNzY3NjU1BiMiJyY1EAAzMhc1IREUDgIjICY1NBMUFjMyNjU0JiMiBnkBQQgdKFZuNyUTDX7A1n1iAQG/xYABBz5wu4/+8uL8g2BnjohoZYNGJzgVHiEWMSNem6y1j9UBCwEarZX8R7y6ajy5jg4Cg6mdoZ6loJ0AAQCSAAAEWQW6ABYAskArDwEfATkBMwIzEEIBQhHeAfkBCQcFFgUkAlgRaBEFAQECExQREhMDFAIBD7gCdEAdAwcJCgoUFQoWAAALCiYICUAgJDSvCQH/CQEJGhi4/8BAFiIkNJAYoBgCcBjwGALvGAEYABQmFhW4/8BADyAkNKAVAfAVARUZFz88GCtOEPRxcis8Tf08ThBdcXIr9nFyKzxN/TwAPzw/PDwQPD/tOTkRFzkDDhA8CDwxMAFdAF0BETYzMh4CFREhETQmJiMiBgYVESERAauIvWGcTx3+5yBRPUZuM/7nBbr95Z9IcIiP/ZECMadaNUSJhv3sBboAAAIAkwAAAawFugADAAcAd7kACf/AQD8RCj9ACVAJAoAJsAnACdAJ7wkFHwlgCX8JoAmwCQUDBgcABQQDDwABQADQAOAAAwBdAgEABgUGBwQKAgcmAQS4/8BACSEkNAQZCD88GCtOEPQrPE39PAA/PD88Pzz9XXE8AwUQPDwQPDwxMAFxXXIrExEhEQERIRGTARn+5wEZBLYBBP78+0oEJvvaAAEAkwAAAawFugADAFO5AAX/wEApEQo/QAVQBQKABbAFwAXQBe8FBR8FYAV/BaAFsAUFAgEAAwAKAgMmAQC4/8BACSEkNAAZBD88GCtOEPQrPE39PAA/PD88MTABcV1yKzMRIRGTARkFuvpGAAEAfgAABpgEPgAnATu5ACn/wEBdEQo/BQYGDBUGFgw0AzQINBg0I0QCRQhFGEQjDCADLylTCWApgCmfKaQGpwemDLUGtQywKdAp4CkOACkvKVApnym/Kd8pBilAGhw0PylQKYAp0CngKQUHIQQHGh0WuAJ0sgoHIbgCdEAeBAcQEREnGxwcJicKAQAGDxAmEhFAWjVgEQFvEQERuAJGQA8aGyYdHEBaNW8cAWAcARy4Aka0JSYmJwG4ASmyAAAnuP/Asw8JPye4/8BANhEKPydAWjUnQEE1J0A8NSdAJCc0J0A6PTQvJ88n3ycDDycfJ4AnAwAnICcwJ/8nBCcZKOM8GCtOEPRdcXIrKysrKysrPE0Q7RD9PPZdcSs8/Tz2cV0rPP08AD88Pzw8EDwQPBA8P+0/7QEREjkAERI5MTABcitxXQBdASsTIRU2MzIWFzY2MzIWFxYVESERNCcmIyIGBhURIRE0JiYjIgYGFREhfgEDi8BmljBGolx1oigd/ucdJ1E7aC7+5x4/NkFoLf7nBCaRqVRVVVRfXESY/VkCX54uPEiLlv4CAkabWixGhJn9/AABAJEAAARZBD4AFgCfQBgHExcTWghoCAS4BAE0CDQQRAhED+kQBQa4AnRAHREHDg0GDAsLAQAKAgEmFgBAICQ0rwAB/wABABoYuP/AQBYiJDSQGKAYAnAY8BgC7xgBGAoLJgwOuAEpsg0NDLj/wEAPICQ0oAwB8AwBDBkXPzwYK04Q9HFyKzxNEO0Q/TxOEF1xciv2cXIrPE39PAA/PDwQPD88P+0xMABdAXFdISERNCYmIyIGBhURIREhFTYzMh4CFQRZ/uckUTlJdCv+5wEFi9Ndmk8fAh6sZThQhLL+HwQmnLRDaIR7AAACAFL/6ASaBD4ADQAZAJdASOgB5wj3E/cVBMcC6AUCEhkFGQkCWRBWE1YWWRiXApgGmAiXDLgJ1QLbBdwJ1QznBecG6A0QpwjLAswGwwjGDAV1CIkGhAgDEbgCdLIKCxe4AnRAFAQHFDkHGmAbcBsCGw4hABkaWEEYK04Q9E3tThBx9k3tAD/tP+0xMABxXQFdcUNYQAlpEGYSZhZpGAQBXVkAXQFdEzQSNjMyABUUACMiJCYlFBYzMjY1NCYjIgZSiv2c8QE0/snskv73igEglm5ulZVubpYCIowBBor+x+/x/sOE/6ieqKignKioAAACAIv+bASXBD4AEAAcAJpALjgTSBMCEjQDOQ05EzQbRANJDUkTRBv5GwlWBlYKWRJWFlYYWRz2B/kbCAEABhq4AnSyBQcUuAJ0QBYLCxAPDhchCBpwHgEeESkODg8mEBABuAEpQAtwAIAAAgAZHT9BGCtOEPRxTe08EP08EOROEHH2Te0APzw/7T/tPzwxMAFdAF0BQ1hADWYGZgppEmYWZhhpHAZdWQBdEyEVNjYzMgAREAAjIiYnESEBFBYzMjY1NCYjIgaLAQYzrmq5AQL+/LlYj0/+5wEWjmZigoZjZ4gEJpxQZP7e/v3+9v7ZRlX96QO5s6uds6einwABAIcAAAM3BD4AEACoQCiXBQEJDgFTBWYFdQUDLxJYDmgOcBIECgkPDB8MAo8M/wwCPwxPDAIMuAJ3QCkHBwEACgMCBgooAAkQCTAJcAkECRp/Ep8SAl8SfxKvEtASBBIQACYBA7gBKUALAgKAAaABAgEZET+5ARwAGCtOEPRxPE0Q7RD9PE4QXXH2XRlN5AAYPzw/PD/tXXFyOTIxMAFdAF1xAEuwF1NLsDVRWlixCjI4WQBdISERIRU2NjMyFwcmIyIGBhEBoP7nAQVDa0RgWVdHPTtSLwQml2tENfUuQar+8QABADD/6AQQBD4AKgLCQMAGEQYjCCcXERcjmBKYFJcnlSoJBxRGFAISuw25Dsch5SP4DfYiBikNVQ1lDZULlxKnIrkMB0EjQCREJmciZCaHEocUhiKDJAk3JkUGRgtKDU8PRiFCIgciJCcmNww1ITUiNSM1JAcGCgURCSEYDScMIiIiIwckIkAscwx4FHkVdil1KogVhCqaFZUqtCK0Iw2AAY8XjBiZKqkqsCwGFyEWQCEjNBZAHB80HxYB3xYBFjMIIVAljyUCJUAYHTQlGiy4/8BAFxEKP1AsATAsAS8sASweITAQARAzASEAuP/Asw8JPwC4/8CzEQo/ALj/wEAJCQ00ABkreLgYK04Q/CsrK03t9HHtThBdcXIr9itxTe30cXIrK+0AsQYCQ1RYQDUGAQEGARYBJiI2IUYhVAFZF2QBaRf2AQoBFwIEGiEiAigTDQwCKBpfBAEERigLUBoBGkYTBz/9XT/9XRESFzkREhc5ERIXOV1xG7kAIv/LsygqNCG4/8uzKCo0Irj/4LMeJDQhuP/gsx8kNCK4/+CzGRo0Ibj/4EAbGRo0aw0BNiJGIpgNlCLEItQiBiEiDA0EBBoAuP/AtRkbNAAzAbj/wLMXLT8BuP+wswkKPgG4/8CzIiU0Abj/wEAdGhw0AAEwAUABUAEEYAGAAfABAwABEAFQAWABBAG4/8CzExY0AbgBAUBNAAQBXwTwBAIERigLFkAZGzQWMxdAFy0/F0AJCj4XQDU3NBdAKy40F0AlKTQXQBocNA8XHxdfF28XBBdVGkAiJDQPGgFQGv8aAhpGEwc//V1xK/RdKysrKysr5Cs//V1x9CtdcXIrKysr5CsREhc5XXErKysrKytZMTABcV0AcXFxcV1dQ1xYuQAk/8lACQsSPw8oCxI/Ibj/7LYNOQwUDDkhuP/ssgw5Irj/6rELOQArKysrASsrWQBxXRMlFhYzMjc2NTQnJickJyY1NDYzMhYXBSYmIyIHBhUUFxYEFxYVFAYjIiYwARoSbmNtNyUUFUn+rFt+2uXa1Cj+9xFfWG8wIBwmAcFZWPTv2f0BLytSVSgcLyAVFBFLPlaZiryOizE+Qh8WIx4VHGZKS4aS0rAAAQAf/+gCkQWdABkAzUApIAAgASMKKQ86DkoOWQ8HGRUAGAMWFQAXEhMUARcSAhQBGAMJBwoHDBi4AQFADwAXoBewFwNgF6AXwBcDF7gBBLIVARS4AnSzABUGB7gCdEAODAsJLwovAAAvAV8BAgG4AQRAKBgDJhcSVRU/FJ8UrxQDYBSAFJAU0BTwFAUAFBAUIBQwFAQUGRp4oBgrThD0XXFyS7A3U0uwO1FaWLkAFP/AOFk8Tfw8/Tz0XTwQ9BnkABg/7T88/TwQ9F1x5BESOREzDw8PDzEwAV0BFSMRFBYWMzI3FwYjIiYmJyY1ESM1MzUlEQJ6wAsnHCdKGGJ8THo5CwmBgQEaBCbg/lSCKxwb2iozUUUxlQHP4NOk/okAAQCN/+gEUwQmABYAnEAXVxFnEZYFAwkGGQY8AjwRSwJLEecCBw+4AnRAEQQLFgAKFRQUCgkGExQmFRUAuAEpQA4WQCAkNK8WAf8WARYaGLj/wEAWIiQ0kBigGAJwGPAYAu8YARgKCyYJCLj/wEAPICQ0oAgB8AgBCBkXPzwYK04Q9HFyKzxN/TxOEF1xciv2cXIrTe08EP08AD88PBA8Pzw/7TEwAF0BXSE1BgYjIiYmNREhERQWFjMyNjY1ESERA046vWlrqkwBGR9SP0hyKgEZn1ViXqqWAqD+GOBlO0915AHA+9oAAAEACwAABFoEJgALARtAFQUoGi80BygaLzQGKBovNAgoGi80A7j/2LMaLzQEuP/AQCAaOjSaBAEGAwsICAoMCxUBFQISAxoJGgoiAC0LxwsMALj/8EAWHSA0CgAFCxQAGQslACoLNAA6C4cACbEGAkNUWLQKAQ0MBLj/wEALCRc0BAEACQEGAAoAPz88ERI5KwEREjk5G0ASCwAKBAsKCQkCAgEGCwAKCTkNuP/AQBgcKDQLDR8NMA1ADQQNFxcaEAo/Ck8KAwq4AjBACwQCOQsEPwRPBAMEugIwAAH/gEAPDDUAASABQAEDARkMxKAYKxlOEPRdKxhN7V3tEP1dGU5FZUTmXSsYTe0APzw/PBA8EDwSOQESOTlZMTABcStdAF0rASsrKysrIQEhExc2NzY3EyEBAbf+VAEnyDoXBg4QygEh/loEJv3itUUWLS0CHvvaAAABAAkAAAY4BCYADAHdQDEACwEKAAYCCgcFCRsAFgIeBBEFGgcUCR4KEQwMEisDKwYjCzkDOQZIA0gGmAOYBgkOuP/AQHcsRzQKAAsEBAUECQsKBAwbABoEFgUUCRkKFQwMIwAoBCcFLQkoCicMMQA3BT4JRgBHAkcFSAdJCXcAeAR3BXgJeAp3DIcAiASHBYgJiAqHDNkA2QTVBdUJ2QrVDOoA6gTkBeQJ6grkDPkA+QT2BfgH9gn5CvYMLbEGAkNUWLQIAQ4NBrj/wLMJITQDuP/AQBUJITQLQAkhNAMLBgMAAQcEAQYJAAoAPzw/PDwREhc5KysrARESOTkbtMILBAUguP9NswYKCSC4/0xAMgMADCALBgMDDAACAQQMAwUKCwcJCAYIBwcFBQQEAgIBBgwKCgkJAAovDj8OAg4XFxoIQQkBDgAgAAYCbQALAm0AQAADAQ60IAEZDcS5ARoAGCtOEPQaGU39Ghj9/RoZ/RhORWVE5l0APzwQPBA8PzwQPBA8EDwQPAEREjk5Ejk5ETk5Ejk5ABEXOSsrK1kxMAFdcSsAXUNcWLQLQA05Brj/+LINOQO4//i2DTkLQAw5Brj/8LIMOQO4//CyDDkGuP/gsgs5A7j/4LELOQArKysrKysrK1kBXQBdIQEhExMhExMhASEDAwFZ/rABEce3AQ+xywEV/qv+8re0BCb9SAK4/UgCuPvaAqv9VQABAA7+UQRSBCYAEwE0tBIoBQETuP/gQBgMDzQIFg0PNAcWDQ80BhYNDzQFFgwPNAK4/8BAHxo6NAUGBgQNCw4GEAIAEwYEEwIEAwMBAQAGE2AQARC4Aa9AEgsPDS8OKAAgFTAVYBUD8BUBFbj/wLMiJjQVuP/AQBIcHjQVFxcaBDkDQBgZNH8DAQO4ASdACQJAGBk0fwIBArgBJ0ASATkAQBw2NCAAMAACABkUxKAYK04Q9F0rTf0Z9F0r9F0rGP1ORWVE5isrcXJNEPTkAD/tXS8/PBA8EDwBEjkROQAREjkSOTkROQcOEDwxMAArASsrKysrXUuwEFNLsDpRWliyBBAAuv/wAAH/8LEDEAE4ODg4WUNcWLkABf/oQA4NET8TEBMZPxMQEhg/Bbj/8LMTGT8FuP/wshIYPwErKysrK1kTIRMTIQEHDgMjIicnFjMyNjcOASv++AEj/olDJUNXf1BRThlCNWJeGQQm/Q4C8vwCuV1iPSIR3A1zWQAAAAABAAAABTXDAAAAAF8PPPUIOQgAAAAAAKLjPB0AAAAA0fjLjfr6/P0QAAgkAAAACQABAAEAAAAAAAEAAAc+/k4AQxAA+vr6ehAAAAEAAAAAAAAAAAAAAAAAAA1dBgABAAAAAAACOQAAAjkAAAKqALgDywBwBHMAEgRzAEYHHQBZBccAWgHnAFwCqgBrAqoAQwMdABwErABVAjkAdQKqAHMCOQCTAjn//QRzAFYEcwCiBHMAMwRzAE0EcwAmBHMAWwRzAFcEcwBXBHMAUwRzAEECqgDJAqoAqgSsAF8ErABVBKwAXwTjAGoHzQA9BccAAAXHAJYFxwBhBccAlAVWAJUE4wCXBjkAYgXHAJYCOQCMBHMAIwXHAJkE4wCdBqoAkQXHAJgGOQBZBVYAlQY5AFkFxwCWBVYASgTjACwFxwCTBVb//weNAAcFVgAABVb//QTjABYCqgCSAjn//QKqACYErABzBHP/7QKqACoEcwBJBOMAhwRzAFUE4wBUBHMAQQKqABgE4wBUBOMAkgI5AJMCOf+iBHMAiQI5AJMHHQB+BOMAkQTjAFIE4wCLBOMAWwMdAIcEcwAwAqoAHwTjAI0EcwALBjkACQRzAAwEcwAOBAAAIgMdADwCPQCwAx0ALQSsAEMFxwAABccAAAXHAGEFVgCVBccAmAY5AFkFxwCTBHMASQRzAEkEcwBJBHMASQRzAEkEcwBJBHMAVQRzAEEEcwBBBHMAQQRzAEECOQCSAjn/6QI5/80COf/QBOMAkQTjAFIE4wBSBOMAUgTjAFIE4wBSBOMAjQTjAI0E4wCNBOMAjQRzAEQDMwBWBHMAVARzAA0EcwA7As0AQgRz//4E4wCLBeX/9wXl//cIAADYAqoAuwKqAAUEZAAxCAD/qgY5AD8FtACYBGQAMgRkADwEZAA8BHMAAQScAG8D9AAsBbQAegaWAKEEZAAAAjEAAAL2ACUC7AAaBiUANwcdAFgE4wBXBOMAZQKqAMMErABVBGQAVARz/+wEZAAfBOUAGgRzAGAEcwBqCAAAyQXHAAAFxwAABjkAWQgAAEgHjQBYBHP//AgAAAAEAACEBAAAaQI5AJgCOQByBGQAMQP0AC8EcwAOBVb/9wFW/qkEc//gAqoASwKqAEsE4wAfBOMAHwRzAEQCOQCTAjkAdQQAAHEIAAABBccAAAVWAJUFxwAABVYAlQVWAJUCOQBqAjn/rgI5/78COf/BBjkAWQY5AFkGOQBZBccAkwXHAJMFxwCTAjkAkwKqAAMCqv/zAqoAEwKqABoCqgDNAqoAkQKqACYCqgBgAqoAOQKqAAME4wAKAjkACgVWAEoEcwAwBOMAFgQAACICPQCwBcf//QTjAFMFVv/3BHMADgVWAJUE4wCLBKwAVQSsAG0CqgBbAqoAGQKqACgGrABcBqwAXAasACgEcwAABjkAYgTjAFQCOQCMBVYASgRzADAFxwBhBHMAVQXHAGEEcwBVBOMAVARr/+0CqgDIBccAAARzAEkFxwAABHMASQXHAJQFwABRBcf//QVWAJUEcwBBBVYAlQRzAEEE4wCdAjkAeQTjAJ0DFQCVBOMAmgPVAJMFxwCYBOMAkQXHAJgE4wCRBjkAWQTjAFIFxwCWAx0AhwXHAJYDHQBQBVYASgRzADAE4wAsAqoAHwTjACwD1QAeBccAkwTjAI0FxwCTBOMAjQTjABYEAAAiBOMAFgQAACIEzwCaBjkAVgaRAFYE6wBOBNoATgPMAE4FeQBOA5IAMAW5AE4Ea//tBNUAuAMrAE8IwAApCAAATwQAAJkIAABPBAAAmQgAAE8EAACYBAAAmAfVAWoFxwCPBKsAVQTVAJ0ErABVBNUCIgTVAQUFq//pBQAByQWrAn4Fq//pBasCfgWr/+kFqwJ+Bav/6QWr/+kFq//pBav/6QWr/+kFqwHABasCfgWrAcAFqwHABav/6QWr/+kFq//pBasCfgWrAcAFqwHABav/6QWr/+kFq//pBasCfgWrAcAFqwHABav/6QWr/+kFq//pBav/6QWr/+kFq//pBav/6QWr/+kFq//pBav/6QWr/+kFq//pBav/6QWr/+kFq//pBav/6QWrAtYFqwBmBav/6gXV//8E1QCSCAAAAAfrATAH6wEgB+sBMAfrASAE1QCyBNUAgATVACoIKwGYCGsBuAdVABAGAAD0BgAAbwRAADoFQAA3BMAAPwQVAEAEAAAlBgAAVQZHAIwEcwCQBav/xwHrAI0D1QCGBxUAIwPpABgE1QCSAtYAXALWAFwE1QCyAtYATQXHAAAEcwBJBccAYQRzAFUFxwBhBHMAVQVWAJUEcwBBBVYAlQRzAEEFVgCVBHMAQQY5AGIE4wBUBjkAYgTjAFQGOQBiBOMAVAXHAJYE4wCSBccABQTjABkCOf+6Ajn/uwI5/9oCOf/aAjn/4QI5/+ICOQBIAjkARwRzACMCOf+iBccAmQRzAIkEcwCNBOMAnQI5/+0FxwCYBOMAkQXJAJwE4wCOBjkAWQTjAFIGOQBZBOMAUgXHAJYDHQAqBVYASgRzADAE4wAsAqoABwXHAJME4wCNBccAkwTjAI0FxwCTBOMAjQXHAJME4wCNB40ABwY5AAkFVv/9BHMADgI5AI0FxwAABHMASQgA/6oHHQBYBjkAPwTjAFcCqgDJB40ABwY5AAkHjQAHBjkACQeNAAcGOQAJBVb//QRzAA4COQCVAqr/1wRzAA0EzQBaBqwAXAasACkGrAAwBqwALwKqALwCqgAmAqoAuwO4//QFx//oBtP/uwc//7sDyv+7Bpn/pgdr/8gGtP+cAjn/KQXHAAAFxwCWBcAAAAVWAJUE4wAWBccAlgI5AIwFxwCZBVYAAAaqAJEFxwCYBSYAZgY5AFkFxwCaBVYAlQTNAFoE4wAsBVb//QVWAAAGeQBWBmoAYgI5/8wFVv//BOsATgOcAE4E4wCOAjkAggSoAGwE4gCQBHMADwOvAE4E4wCOBFMATgI5AJMEdgCOBHMADwTlAJAEcwALA5AATgTjAFIE8wB2BCkATgSoAHYEmwARBgcAdgbCAE4COf/NBKgAdgTjAE4EqAB2BsIATgVaAJcHFQAvBIkApAWxAFgFVgBKAjkAjAI1/8oEcwAjCMAAGgiAAJ0HAAA3BOIAmgT6AAAFwACZBccAAAXAAJsFxwCWBIkApAWz//oFVgCVBzsAFwUDACwFwACZBcAAmQTiAJoFnQAgBqoAkQXHAJYGOQBZBcAAmQVWAJUFxwBhBOMALAT6AAAG1ABZBVYAAAXYAJoFnwB9CAoAmggnAJoG9QAaB9UAnQXAAJsFsQBXCEAAlgXAAAQEcwBJBPEAXATrAJYDVQCIBRT/+QRzAEEFrP//A/oAGATrAIwE6wCMBAEAiAUVABkF6wCbBNUAiATjAFIE1QCIBOMAiwRzAFUD6wAVBHMADgcAAFQEcwAMBOsAiQSlAHIGqwCMBsAAjQXVACgG1QCVBOsAmQRrADgG1QCRBKv/+wRzAEUE4wAAA1UAiARrAFEEcwAwAjkAkwJA/9ACOf+iB8AAGAdAAIwE4wAABAEAiARzABIE1QCIA+UAlgOTAIgIAABBCOsAowYgADAAAAEBAAAAHgAAADEAAAAxAAABAQAAAH8AAAB+AAAAjAAAAIwAAAEBAAAAEAAAAQEAAAEhA5MAfQAAAIwCZQDIAAADAgAA/wECqgDJBKkAWQSbAEEDpwAKBGYAMgTqAIICLwCHA04AWgTtAIcFAwB9Ai8AhwQsACgD7QBLA/gAQQTjAIcFCgA3Ai8AhwMWAEsE6ABQBFkACgTAAGQEsgBkA/8ACgQYAAoElQCCBCwAKAW4AFoFYwAtBF4AhwReAIcEXgCHAjYAUAQJAFAGiwCHAi//rAQsACgELAAoA/j/FgP4/xYEeQAyBbgAWgW4AFoFuABaBbgAWgSpAFkEqQBZBKkAWQSbAEEDogAKBGYAMgTqAIIClQAAA4EAAAUDAH0ClQAABCwAKAPtAEsD+ABBBQoANwMWAEsE6ABQBMAAZASyAGQEGAAKBJUAggQsACgFuABaBWMALQIvAIcEmwBBA+0ASwSyAGQE2wBBAAD/3AAA/yUAAP/cAAD+UQKNAKsCjQCgAtoAQwPAAH4Blv+6AAAARgAAAEYAAABGAAAARgAAAEgAAABGAAAARgAAAEYEfgGIBH4BUAR+AQQEfgCeBH4BLQR+AOoEfgDVBH4AnAR+ALwEfgDuBDUAhQKNAMEENQCzBgABAAYAAQACvgBYBgABAAR+AKUEfgC9BH4A3gYAAQAGAAEABgABAAYAAQAGAAEAAAAARgYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABOb/ugYAAQAGAAEABgABAAUyADkFMgA5Aiz/ugIs/7oGAAEABgABAAYAAQAGAAEABJ4ANAR4ADAEMP+6BDD/ugN2AAoDdgAKBg4AKQcIACkC4v+6BFb/ugYOACkHCAApAuL/ugRW/7oFKACXBG8ACgNSAAMGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAAAAAwAAAARgAAAEYAAABAAAAARgYAAQAGAAEAAAD/3AAA/lEAAP8WAAD/FgAA/xYAAP8WAAD/FgAA/xYAAP8WAAD/FgAA/xYAAP/cAAD/FgAA/9wAAP8gAAD/3ARzAC0IAAAABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAKNAH8CjQBnBgABAAWgAC4DwAB+AegAAAIH/8MBvABeAeD/+gOcAAYDnAAGAbwAXgHgABoFKACXBJ4AEQIs/7oCLP+6AbwAiAHgABoFMgA5BTIAOQIs/7oCLP+6Ar4ANgNSAAMFMgA5BTIAOQIs/7oCLP+6BTIAPAUyADwCLP+6Aiz/ugSeADQEeAAwBDD/ugQw/7oEngA0BHgAMAQw/7oEMP+6BJ4ANAR4ADAEMP+6BDD/ugK+AGkCvgBpAr4AaQK+AGkDdgAKA3YACgN2AAoDdgAKBzIAQAcyAEAE3v+6BN7/ugcyAEAHMgBABN7/ugTe/7oIgABACIAAQAYs/7oGLP+6CIAAQAiAAEAGLP+6Biz/ugQw/7oEMP+6BDD/ugQw/7oEMP+6BDD/ugQw/7oEMP+6BFQANAPAAEYEVP+6AuL/ugRUADQDwABGBFT/ugLi/7oGEAAvBhAALwJw/7oCmP+6BOYAJwTmACcCcP+6Apj/ugRUACkEVAApAuL/ugLi/7oDnAAjA5wAIwHg/7oB4P+6AuIAIQLiACEDUv+6A1L/ugRUAD4EVAA+Aiz/ugIs/7oCvgBYA1IAAwPA/7oDnP+6A5wABgOcAAYFKACXBG8ACgUoAJcEngARAiz/ugIs/7oEVAAABMQAAAPkACIEVAAaA+QAIgRUABoD5AAiBFQAGgYAAQAGAAEAAAAARgAAAEYGAAEABgABAAYAAQAAAABGAAAARgYAAQAGAAEAAAAASAAAAEYGAAEABgABAAYAAQAAAABGAAAARgAAAEYAAABGAAAAQAAAADAGAAEAAAAARgAAAEYGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQACjQDKAo0AxwKNAMYGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAK+AGkBAP+6CAD/uhAA/7sG0wBZBbAAUgajAJMFywCNAAD9iAAA+8EAAPxfAAD+MQAA/K0AAP1VAAD+JgAA/fEAAP0YAAD8aQAA/ZUAAPvgAAD8cAAA/tQAAP7NAAD+oAQbAHgGrABcBqwAGQAA/kUAAP1VAAD9pgAA/F8AAP4lAAD9GAAA++AAAPr6AAD7NgAA/HAAAPuHAAD7mwAA/M4AAPxUAAD7wwAA/JQAAPv1AAD9sAAA/lkAAP1+AAD8ggAA/TQAAP5QAAD+RgAA/NEAAP0+AAD9AgAA/DoAAPzpAAD8JgAA/AcAAPwvAAD7ngAA+3YCOQCTBccAAARzAEkFxwAABHMASQXHAAAEcwBJBccAAARzAEkFxwAABHMASQXHAAAEcwBJBccAAARzAEkFxwAABHMASQXHAAAEcwBJBccAAARzAEkFxwAABHMASQXHAAAEcwBJBVYAlQRzAEEFVgCVBHMAQQVWAJUEcwBBBVYAlQRzAEEFVgCVBHMAQQVWAJUEcwBBBVYAlQRzAEEFVgCVBHMAQQI5AGoCOQBdAjkAjAI5AJMGOQBZBOMAUgY5AFkE4wBSBjkAWQTjAFIGOQBZBOMAUgY5AFkE4wBSBjkAWQTjAFIGOQBZBOMAUgbTAFkFsABSBtMAWQWwAFIG0wBZBbAAUgbTAFkFsABSBtMAWQWwAFIFxwCTBOMAjQXHAJME4wCNBqMAkwXLAI0GowCTBcsAjQajAJMFywCNBqMAkwXLAI0GowCTBcsAjQVW//0EcwAOBVb//QRzAA4FVv/9BHMADgXHAAAEcwBJAjn/ygI5/8oGOQBZBOMAUgXHAJME4wCNBccAkwTjAI0FxwCTBOMAjQXHAJME4wCNBccAkwTjAI0AAP75AAD++QAA/vQAAP7vBIn//QNVAAcHOwAXBaz//wTiAJoEAQCIBOIAmgQBAIgFxwCWBNUAiARzAAEEcwASBHMAAQRzABIFVgAABHMADAWfAH0EpQByBZ8AnATjAJIFzwBZBHMATAY5AFYE4wBSBTIAOQIs/7oCcP+6Apj/ugTmACcCLABlAiwAFgIsABYCLAARAiwAQwIs/9IAAP7wAAAADwAA//UCqgCQAqoAkAAAAAAAAABeAAAAXgAA/8sBvAAPAeD/vwG8//UB4P/NAbwAHQHgAAkBvACIAeAAGgOcAAYDnAAGA5wABgOcAAYFKACXBG8ACgUyADkFMgA5Aiz/ugIs/7oFMgA5BTIAOQIs/7oCLP+6BTIAOQUyADkCLP+6Aiz/ugUyADkFMgA5Aiz/ugIs/7oFMgA5BTIAOQIs/7oCLP+6BTIAOQUyADkCLP+6Aiz/ugUyADkFMgA5Aiz/ugIs/7oEngA0BHgAMAQw/7oEMP+6BJ4ANAR4ADAEMP+6BDD/ugSeADQEeAAwBDD/ugQw/7oEngA0BHgAMAQw/7oEMP+6BJ4ANAR4ADAEMP+6BDD/ugSeADQEeAAwBDD/ugQw/7oCvgBPAr4ATwK+AGkCvgBpAr4AaQK+AGkCvgBPAr4ATwK+AGYCvgBmAr4AaQK+AGkCvgBpAr4AaQK+AC8CvgAvAr4AIgK+ACIDdgAKA3YACgN2AAoDdgAKA3YACgN2AAoDdgAKA3YACgN2AAoDdgAKA3YACgN2AAoDdgAKA3YACgN2AAoDdgAKBzIAQAcyAEAE3v+6BN7/ugcyAEAHMgBABN7/ugTe/7oHMgBABzIAQATe/7oE3v+6CIAAQAiAAEAGLP+6Biz/ugiAAEAIgABABiz/ugYs/7oEMP+6BDD/ugRUADQDwABGBFT/ugLi/7oGEAAvBhAALwYQAC8CcP+6Apj/ugYQAC8GEAAvAnD/ugKY/7oGEAAvBhAALwJw/7oCmP+6BhAALwYQAC8CcP+6Apj/ugYQAC8GEAAvAnD/ugKY/7oE5gAnBOYAJwTmACcE5gAnCT4AMgk+ADIHQP+6B0D/ugYOACkHCAApAuL/ugRW/7oEVAApBFQAKQLi/7oC4v+6BFQAKQRUACkC4v+6AuL/ugRUACkEVAApAuL/ugLi/7oGDgApBwgAKQLi/7oEVv+6Bg4AKQcIACkC4v+6BFb/ugYOACkHCAApAuL/ugRW/7oGDgApBwgAKQLi/7oEVv+6Bg4AKQcIACkC4v+6BFb/ugOcACMDnAAjAeD/ugHg/7oDnAAjA5wAIwHg/7EB4P+xA5wAIwOcACMB4P+6AeD/ugOcACMDnAAjAeD/ugHg/7oEVAA+BFQAPgIs/7oCLP+6BFQAPgRUAD4EVAA+BFQAPgRUAD4EVAA+Aiz/ugIs/7oEVAA+BFQAPgSeADQEeAAwBDD/ugQw/7oCvgBYA1IAAwMaABoDGgAaAxoAGgOcAAYDnAAGA5wABgOcAAYDnAAGA5wABgOcAAYDnAAGA5wABgOcAAYDnAAGA5wABgOcAAYDnAAGA5wABgOcAAYFKABCBG//2QUoAJcEbwAKAiz/ugIs/7oDnAAGA5wABgUoAJcEbwAKAiz/ugIs/7oFKACXBG8ACgZ/AEQGfwBFBn8ARAZ/AEUBqAAoAAD+KQAA/owAAP8lAAD/IwAA/voAAP96AAD+WQj8ADIIrQAyAAD/tQAA/7YAAP7wAAD/WQAA/lkAAP+MAbQAAAL3AAAAAP6FAAD/BwTNADIAAP9YAAD/WAAA/1kHMgBABzIAQATe/7oE3v+6CIAAQAiAAEAGLP+6Biz/ugRUADQDwABGBFT/ugLi/7oDwAB+AuIAIQK+AFgCLP+6ApD/ugH0AC8B9AA7AfQAEgH0ALEB9ABtBg4AKQcIACkCLwCHAAD+yANQAAAEXgCHA+T/9QRU//UD5AAiBFQAGgPkACIEVAAaA+QAIgRUABoD5AAiBFQAGgPkACIEVAAaA+QAIgRUABoEfgByBH4AvQPkAA8EVAAPBOMAGwaxAB4FwACbBOMAhwXAAAoE4wAKBccAaQXHAGEEcwBVBcf//QazAB4FwABcBOMAVATaAE4FVgBmBQMAbwTj/6wGOQBiBRgAAgdyAJICOQCTAjkABwXHAJkEcwCJAjkAGwRzAA8H7wCWBcf/rQTjAI4GOQBWBxgAWQXzAFUGQQAeBOMAiwVWAJUFVgBkBHMAYwTNAFoC4QAeAqoAHwTjABgCqgAfBOMALQZqAGIFxwCTBikAAARzAA4E4wAWBAAAIgTjADoE4wBZBDYAKgQ2ADkEcwAzBHMAWwP6AB4EogAfBOMAiwI9ALAD+wCwBK0AVgKqALgKqgCUCccAlAjjAFQJVgCdBxwAnQRyAJMKOgCYCAAAmAccAJEEcwBMBccAAARzAEkAAP7+BccAAARzAEkIAP+qBx0AWAY5AGIE4wAkBjkAYgTjAFQFxwCZBHMAiQY5AFkE4wBSBjkAWQTjAFIE4wA6BDYAIgI5/6IKqgCUCccAlAjjAFQGOQBiBOMAVAhDAJYFUgCVBccAmATjAJEFxwAABHMASQXHAAAEcwBJBVYAlQRzAEEFVgCVBHMAQQI5/zcCOf8tAjn/9AI5/+YGOQBZBOMAUgY5AFkE4wBSBccAlgMd/80FxwCWAx0AgAXHAJME4wBnBccAkwTjAI0FVgBKBHMAMATjACwCqgAfBJ4ALgQpAEkFxwCWBOMAkgWfAJwFDABSBQwAUgTjABYEAAAiBccAAARzAEkFVgCVBHMAQQY5AFkE4wBSAAD+/QY5AFkE4wBSBjkAWQTjAFIGOQBZBOMAUgVW//0EcwAOBHMARQTjAFQE4wCCBOMAhwRzADQEcwAUBOMAVATjAFQEcwBMBkEATAP6AE8D+gAYBYcAGASKAFICqv/EBOMAVATjAFQEsABSBHMADwTOAA8E4wCKBOMAkgTjAJICOQAbAjkAawM+AEQCqAAAAtkAFAI5AJME1ACTBx0AhQcdAIUHHQB+BOP/pgTjAJEE6wCMBOMAUgarAFIGwgBOBf8AUgMd/+YDHf/mAx3/5gMdAIcDHQCHAx0AhwMd/+YEqwCKBKsAigRzADACqv/EAqr/xAKq/5sEUQAeAqoAGQKqAB8E4wAbBPgASwSoAJEEcwASBjkACQRzAA8EkQAPBAAAIgVwACIENgAiBDYAIgRzAEIEcwBVBHMAQgRzAFUGOQBZBOsAlgSKAE8EsABSBNUAiAOrAB4EcwAUA54AiATjAFsEcwBCBHMAVQg/AFQHiQBUCa8AVAaCAB8ERgAfBpgAHwb0ABgGNQCTBYoAkwRFAB4EggCIAvEAMgLxADIBjv/iAgQAMgIEAAACBAAAAwAAMgQvAAAC4gAAAecAXAPLAHACOQCYAjkAdQI5AJQCqgDzAqoA8wMAADIDAAAyBKwAXwSsAF8ErAAqBKwAKgKqASECqgC7AqoAKgKqASECqgATAqoAKgKqALsCqgDKAqoAygKqAPMCqgDzAqoApgKqAKYCqgCmAqoAEwKq/+ECqv/7Au0AAAEhADIDAgAyAu4AAAMAADIDEACWAxAAlgMQAJYDEACWAxAAlgKqAGICqgBiAqoAAwKqAB0EAABpBFcAlgRXAJYEVwCWBFcAlgRXAEMEVwBDBFcAQwRXAEMEVwBDAxAAQwRXAC8EVwAvBFcALwRXAC8EVwAvAxAALwRXACUEVwAlBFcAJQRXACUEVwAlAxAALwRXABoEVwAaBFcAGgRXABoEVwAaAxAAGgRXAEIEVwBCBFcAQgRXAEIEVwBCAxAAQgRXAJYEVwCWBFcAlgRXAJYEVwBCBFcAQgRXAEIEVwBCBFcAQgMQAEIEVwAvBFcALwRXAC8EVwAvBFcALwMQAC8EVwAvBFcALwRXAC8EVwAvBFcALwMQAC8EVwAmBFcAJgRXACYEVwAmBFcAJgMQACYEVwBCBFcAQgRXAEIEVwBCBFcAQgMQAEIEVwCWBFcAlgRXAJYEVwCWBFcAQgRXAEIEVwBCBFcAQgRXAEIDEABCBFcAJgRXACYEVwAmBFcAJgRXACYDEAAmBFcAIwRXACMEVwAjBFcAIwRXACMDEAAjBFcALwRXAC8EVwAvBFcALwRXAC8DEAAvBFcASwRXAEsEVwBLBFcASwRXAEsDEABLBFcAlgRXAJYEVwCWBFcAlgRXAEIEVwBCBFcAQgRXAEIEVwBCAxAAQgRXABoEVwAaBFcAGgRXABoEVwAaAxAAGgRXACQEVwAkBFcAJARXACQEVwAkAxAAJARXAC8EVwAvBFcALwRXAC8EVwAvAxAALwRXAE4EVwBOBFcATgRXAE4EVwBOAxAATgRXAJYEVwCWBFcAlgRXAJYAAP6vAAD+vwAA/bUAAP7IAAD/eAAA/rEAAP89AAD+bwAA/q4AAP/OAAD/ZgAA/m8AAP7IAAD+yAAA/2gAAP9oAAD/aAAAAAAAAP8fAAD/HwAA/0QAAP9fAAD+hwAA/+wAAP+cAAD/UQAA/1EAAP9RAAD+vwAA/xUAAAAAAAD+sQAA/z0AAP9rAAD+8gAA/0cAAP/OAAD+hwAA/rsAAP6uAAD+rgAA/sgAAP7IAAD+pgAA/r8AAP23AAD+vgAA/qYAAP6/AAD9tQAA/h8AAP7iAAD/nAAA/ocAAP9EAAD+ugAA/yMAAP+aAAD9uQAA/jsAAAAAAAD+pwAA/2gAAP4XAAD/dAAA/ocAAP4AAAD/ZgAA/0QAAP6nAAD+pwAA/qcAAP8DAAD/UgAA/R8AAP9TAAD/UwAA/1MAAP6xAAD+sAAA/6EAAP6MAAD+uAAA/q8AAP6iAAD+ugAA/fQAAP8ZAAD/LQAA/owAAP6IAqoAuwKqACoCqgDIBOIAZwSoAAoGKQAACAIAAAYpAAAF/wBSBsIATgVpABQGOQBZBOMAUgXHAHcEcwBVBOMAlwOeAIgGAwAABDwAHQZvAAoE4gAKB+8AlgcdAIUFnwB9BOMAigWfAJwE1wAKBVYAZAVWAGQFJAAUBNQACgXhAFUEoABLBA4AFAOEACgFaQAUBPEAXARzAFUCOf+iBjkAVgPUAFED1ABRBVYAlQXAAJkEcwBBBOsAjAo9AFkGOgAUBvQAGgWfABsHzgCMBl4AkwVWAAAEcwALB2gAjAZnAJMGeQBWBgcAdgieAIwH2ACTBQMARgP6AEMGeQBWBgcAdgY5AFYE4wBSBoX//wUsAAsGhf//BSwACwj2AFkHywBSBoQAIwUaACMKPQBZBzUAVQAA/jcKPQBZBjoAFAXHAGEEcwBVBKwADwAA/qYAAP6xAAD/jQAA/40AAPwrAAD8TAXAAJkE6wCMBcAAEQTrABsFVgCVBOMAiwWfAJwEyQCIBQMALAP6ABgE4gARBAEADQYXABoE/AAoBwkAlgW2AIgJAgCZB18AiAXHADsEnwA0BccAYQRzAFUE4wAtA+sAFQbSACwFgwAVBZ8AfQSlAHIG2gAKBW0ACgbaAAoFbQAKAjkAjAc7ABcFrP//BZ0AmgTIAIgFnQAgBRUAGQXHAJYE1QCIBccAlgTVAIgFnwB9BKUAcgaqAJEF6wCbAqoAGgXHAAAEcwBJBccAAARzAEkIAP+qBx0AWAVWAJUEcwBBBc8AWQRzAEwHOwAXBaz//wUDACwD+gAYBQMALAQ2ACIFwACZBOsAjAXAAJkE6wCMBjkAWQTjAFIGOQBWBOMAUgWxAFcEawA4BPoAAARzAA4E+gAABHMADgT6AAAEcwAOBZ8AfQSlAHIH1QCdBtUAlQXAAF4E4wBUCD4AXgd6AFQHrQBGBsQAQwVDAEYESgBDCBoAIAelABkIQwCWB2YAiAY5AGIEsABSBiAALQWbABUAAP9DAAD+yQAA/3cAAP+wAAD/RwAA/1YAAP90AAD+1wAA/qwAAAAAAAD/UgAA/1YAAAAAAAD+rAAA/ZoAAAAAAAD/agAA/3wAAP9pAAD/VgAA/qwAAP9/AAD/VgAA/e8AAP9DAAD/aQAA/3wAAAAAAAD9rgAA/4wAAAECAAD+7wAA/u8AAP79AAD++QAA/1MAAP74AAD++QXHAAAEcwBJBccAlgTjAIcFxwCWBOMAhwXHAJYE4wCHBccAYQRzAFUFxwCUBOMAVAXHAJQE4wBUBccAlATjAFQFxwCUBOMAVAXHAJQE4wBUBVYAlQRzAEEFVgCVBHMAQQVWAJUEcwBBBVYAlQRzAEEFVgCVBHMAQQTjAJcCqgAYBjkAYgTjAFQFxwCWBOMAkgXHAJYE4wCSBccAlgTjAJIFxwBOBOMAOwXHAJYE4wCSAjn/0gI5/9ICOQAbAjn/zgXHAJkEcwCJBccAmQRzAIkFxwCZBHMAiQTjAJ0COQCTBOMAnQI5/+sE4wCdAjn/3QTjAJ0COf/LBqoAkQcdAH4GqgCRBx0AfgaqAJEHHQB+BccAmATjAJEFxwCYBOMAkQXHAJgE4wCRBccAmATjAJEGOQBZBOMAUgY5AFkE4wBSBjkAWQTjAFIGOQBZBOMAUgVWAJUE4wCLBVYAlQTjAIsFxwCWAx0AhwXHAJYDHQCHBccAlgMdAIcFxwCWAx0AWQVWAEoEcwAwBVYASgRzADAFVgBKBHMAMAVWAEoEcwAwBVYASgRzADAE4wAsAqoAHwTjACwCqgAfBOMALAKqAB8E4wAsAqoAHwXHAJME4wCNBccAkwTjAI0FxwCTBOMAjQXHAJME4wCNBccAkwTjAI0FVv//BHMACwVW//8EcwALB40ABwY5AAkHjQAHBjkACQVWAAAEcwAMBVYAAARzAAwFVv/9BHMADgTjABYEAAAiBOMAFgQAACIE4wAWBAAAIgTjAJICqv/eBjkACQRzAA4EcwBJAjkAjQTrAE4E6wBOBOsATgTrAE4E6wBOBOsATgTrAE4E6wBOBccAAAXHAAAG8//yBvMAAAbz//IG8wAABvMAQwbzAEMDzABOA8wATgPMAE4DzABOA8wATgPMAE4GHv/yBh4AAAeu//IHrgAAB67/8geuAAAE4wCOBOMAjgTjAI4E4wCOBOMAjgTjAI4E4wCOBOMAjgaP//IGjwAACB//8ggfAAAIH//yCB8AAAgfABQIHwAUAjkAkAI5AJACOf+2Ajn/xAI5/94COf/sAjn/swI5/8ADAf/yAwEAAASR//IEkQAABJH/8gSRAAAEkQAUBJEAFATjAFIE4wBSBOMAUgTjAFIE4wBSBOMAUgad//IGnQAACFX/8ghVAAAHyf/yB8kAAASoAHYEqAB2BKgAdgSoAHYEqAB2BKgAdgSoAHYEqAB2BoIAAAf+AAAIYgAAB67/8wbCAE4GwgBOBsIATgbCAE4GwgBOBsIATgbCAE4GwgBOBs7/8gbOAAAIhv/yCIYAAAf6//IH+gAAB/r/8wf6//ME6wBOBOsATgPMAE4DzABOBOMAjgTjAI4COf/nAjkAjQTjAFIE4wBSBKgAdgSoAHYGwgBOBsIATgTrAE4E6wBOBOsATgTrAE4E6wBOBOsATgTrAE4E6wBOBccAAAXHAAAG8//yBvMAAAbz//IG8wAABvMAQwbzAEME4wCMBOMAjATjAIwE4wCMBOMAjATjAIwE4wCMBOMAjAaP//IGjwAACB//8ggfAAAIH//yCB8AAAgf//MIH//zBsIATgbCAE4GwgBOBsIATgbCAE4GwgBOBsIATgbCAE4Gzv/yBs4AAAiG//IIhgAAB/r/8gf6AAAH+v/zB/r/8wTrAE4E6wBOBOsATgTrAE4E6wBOBOsATgTrAE4FxwAABccAAAXH/9EFx//dBccAAAKqANwCqgDKAqoA3AKq//MCqv/zBOMAjATjAIwE4wCMBOMAjgTjAIwG5gAABuYAAAdXAAAHVwAABccAlgKq//ICqv/yAqr/8wI5/+UCOf/bAjn/zgI5/84COf/CAjn/uwI5/+gCOf/eA8kAAAPJAAACqgAAAqoAAAKq//MEqAB2BKgAdgSoAHYEqAB2BPMAdgTzAHYEqAB2BKgAdgVW//0FVv/9Bub/2AdK/90GHgAAA7j/9AO4//QCqgAqBsIATgbCAE4GwgBOBsIATgbCAE4HZf/RBp3/3QeW/9EGzv/dBmoAYgKqALsCqgDcBHMACgXHAGEFxwBhBx0AfgXHACEJzQCWB40ABwXHACAE4wAtCLAAFAQAADAEwQBmAAD/UwAA/1MAAP9TAAD/UwI5ABsCOf+iBHMAAAVWABIGswBUA/4AVwarAJEEDAAfBdb/5gXW/+YCqgCEAqoAhAKqAMkCqgDJAqoAkQKqACoCqv/FAqr/wwKq//MCqgDJAqoAqQKqAKkCqgCpAqoAqQMuAB4DLgAeAqoAOgAA/3MAAP+dAAD+yAAA/yMAAP9yAAD/cgAA/ucAAP+dAAD/UwAA/1MAAP9TBVYAlQTjAIsEtQAABjUAAAcdAGEE6wAPBHMAVQSZAJEEmQAbBAEAjAP6ABgCOQCTBA8ASQR2AI4DngAOBesAmwTrAIwE4wBSBHMANATxAFIE8QBSBPEAIQeNAFQEkgBLBOMAUwTjAFME6QCMBKv/+wSr//sD6wAVBKgAdgTjAFEGJABRBOAAUQRzAAsGOQAJBAAAIgPfACID8gBLBOwAFANVAIgEcwASBNUAiATpAIwGBwB2BRUAGQPjAAAFkQAAA6IAMgOiAAADowAyA1UAMgNVADIEAwAyA3wAMgFyAFUC3gAyA7AAMgMeADIEIgAyA3cAMgN4ADIEJgAyA3oAMgNbADIDrAAyA3cAMgN7ADIFFAAAAwUAMgMFADIDIQAyBLYAMgMhADIDIQAyAwIAMgMCADICzwAyAs8AMgMgADIBIQAyAsoAMgSEADQC8gAyA0gAMgMKADIDSQAyA0kAMgMgADIBvAAKAvIAMgNCADIEhAAyAukAAANMAAoDGwAyAukAAANDADID2gAyAwgAAAEhADICBAAyAvIAMgLpAAADGwAyAukAAANCADID2gAyAwgAAAXtAEYKmABGBhMARgaJ/7oFQf+6AekAHgRUABAAAP8NAAD/NQAA/s4AAP63AAD+yQAA/8cAAP9PAAD/ngAA/vACvgBpAr4AaQN2AAoDdgAKA8D/ugOc/7oDwP+6A5z/ugXIADkFkgAyBhYAggUZAEsFJABBBg8AhwVYACgGjwAtBKwAVQAA/jsAAP5mAAD+aARz//wEAACEA9X/ugHg/7oB4P+xAeD/ugHg/7oG0AAuCYQAIwQAAAAIAAAABAAAAAgAAAACqwAAAgAAAAFVAAAEcwAAAjkAAAGaAAAAqwAAAAAAAAXl//cFxwBhBqoAkQXrAJsHYACNB6EAVAehAFsFxwAABccAYQRzABQE4wARBOMALARzADkEAAAiBSkAQgAAAQEAAP9CAAD+rQAA/zoAAP9TBPMACgXHAGkFxwBhBccAaQSJAKQDVQCIAAD/QwAA/wEAAP+sAxYAfQAA/zcCmP+6Az0AHgAA/zoAAP9IAAD/SQAA/34AAP9PAAD/SgAA/p4FMgA5BTIAOQIs/7YCLP+2BTIAPAUyADwCLP+6Aiz/ugUyADkFMgA5Aiz/ugIs/7oFMgA5BTIAOQIs/7oCLP+6BTIAOQUyADkCLP+6Aiz/ugUyADkFMgA5Aiz/ugIs/7oFMgA5BTIAOQIs/7oCLP+6BJ4ANAR4ADAEMP+6BDD/ugSeADQEeAAwBDD/ugQw/7oCvgBPAr4ATwK+AGkCvgBpA3YACgN2AAoHMgBABzIAQATe/7oE3v+6BFQANAPAAEYEVP+6AuL/ugRUADQDwABGBFT/ugLi/7oEVAA0A8AARgRU/7oC4v+6BhAALwYQAC8CcP+6Apj/ugYQAC8GEAAvAnD/ugKY/7oGDgApBwgAKQLi/7oEVv+6Bg4AKQcIACkC4v+6BFb/ugYOACkHCAApAuL/ugRW/7oC4gAhAuIAIQNS/7oDUv+6AuIAIQLiACEDUv+6A1L/ugRUAD4EVAA+Aiz/ugIs/7oEVAA+BFQAPgIs/7oCLP+6BFQAPgRUAD4CLP+6Aiz/ugOcACMDnAAjAeD/ugHg/7oDdgAKA3YACgN2AAoDdgAKBzIAQAcyAEAE3v+6BN7/ugTj/8EE4wBUAqr/8wcd/8EE4//VBOP/xQMd/8EDHf/BBHP//wKq/9oEAAAhBOMAgwLwADIE3ABOBvsAHwI5ABsCOQAbBOMAFASoABQE+AAUBOMAhwTjAFQCqgAYBiUAVARzAIkCOQBwBx0AfgTjAJEE4wCLAx0AZgRzADADuv/EBHMACwRzAAwEAAAiBHMASQTjAFQE4wBUBHMAQQP6AE8D+gAYBT4AUQI5AJMEcwA0Aqr/xATjAI0ENgAiAyEAMgMKADIDCgAGA0gAMgLPADIB8AAKAfAAAAMgADIC8QAyAXQACgEhADIBIQAyAXQACgJ2AAABjgAyAVAAMgJJADIEhAA0BIQAMgNfAAADXwAyAvoAMgNIADIEAwAyAwIAMgI5AAABvAAKA0AACgNeADIC6gAyAuoAMgLpAAAC5AAyAuQAMgO+ADIDCgAyAugAMgAA/pIAAP6SAAD/cwAA/p8CqgDJAwUAMgMCADIDSAAyAu4AAAMCADIGOQBiBccAAAVWAB4FxwBhAqoAQQTrAE4E6wBOBOsATgTrAE4E6wBOBOsATgTrAE4E6wBOAjn/tgI5/7YCOf/EAjn/xAI5/7YCOf+2Ajn/xAI5/8QEqAB2BKgAdgSoAHYEqAB2BKgAdgSoAHYEqAB2BKgAdgI5/8kCOf/JAjn/yQI5/8kEqAB2BKgAdgSoAHYEqAB2A+QAIgRUABoD3wAwBcf//QXHABYFVgAABVYAlQRzAEEEcwAjAjn/ogYzAFkE4wBbBccAAAMdABsFVv/9BHMADgRzADQEcwBVBHMANAI5AJMEiQARA1UAGwVWAAAEcwAMBVYAAARzAAwFAwBvA/oATwWdACAFFQAZAAD+xgAA/tQAAP7GAAD+1AAA/l8AAP5fAAD/cgAA/3MAAP7nCAAAAAQBAF0EcwA0BOMAEQI5ABsE4wAGBVb//QXHAJYEcwBJAqr/zQXHAJYE4wCSBccAmQRzAIkE4wAWBAAAIgRzACgEVACWA3wAiAW5AE4AAP9TAAD/vAAA/v4AAP7+AAD+pAAA/qQCOQCTBckAnAXHAJgFyQCcAAD+4AAA/zAAAP7UAAD+1QAA/sAAAP7QAAD+2AAA/tgAAP7YAAD+2AAA/cYGOQBZBOMAWweNAAcGOQAJBbkAkQAA/psGGwBZBNkABghbAAcG3gAGAqoAyQMcAFUB5wBcAecAXAQAAJkEAACZAqoAuAKqALgCqgC4AqoAAwTjACwEcwArBMMACgRzABQGlwCHBzgAUAAAAAAAAABsAAAAbAAAAGwAAABsAAAAbAAAAGwAAABsAAAAbAAAAGwAAABsAAAAbAAAAGwAAABsAAAAbAAAAGwAAABsAAAAbAAAAKoAAAEAAAACBAAAAoYAAAQsAAAFhAAABp4AAAgQAAAJRAAACgAAAAueAAAM5AAADOQAAAzkAAAM5AAADOQAAAzkAAAM5AAADOQAAA5eAAAPxgAAEQAAABHqAAASqAAAE0QAABSKAAAVXgAAFeYAABaEAAAYTgAAGKoAABr+AAAc/AAAHgQAAB7UAAAe1AAAIDgAACKYAAAjLgAAJA4AACQOAAAkDgAAJA4AACUEAAAlBAAAJXgAACV4AAAleAAAJXgAACV4AAAleAAAJ4YAACiCAAApvgAAKq4AACy6AAAtugAAL5YAADCWAAAxOAAAMTgAADE4AAAxpAAAM1gAADRCAAA1MgAANi4AADYuAAA3EgAAOlgAADt4AAA8YAAAPbQAAD/QAAA/0AAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAABBTgAAQU4AAEFOAAEAAA1dAPIAPACPAAYAAgAQAC8AVQAABzz//wAFAAIAAAAUAPYAAQAAAAAAAAAQAAAAAQAAAAAAAQARABAAAQAAAAAAAgAHACEAAQAAAAAAAwARACgAAQAAAAAABAARADkAAQAAAAAABQAMAEoAAQAAAAAABgARAFYAAQAAAAAABwAHAGcAAQAAAAAACAAHAG4AAQAAAAAACQAHAHUAAwABBAkAAAAgAHwAAwABBAkAAQAiAJwAAwABBAkAAgAOAL4AAwABBAkAAwAiAMwAAwABBAkABAAiAO4AAwABBAkABQAYARAAAwABBAkABgAiASgAAwABBAkABwAOAUoAAwABBAkACAAOAVgAAwABBAkACQAOAWZPcmlnaW5hbCBsaWNlbmNlQkVGTkhDK0FyaWFsLEJvbGRVbmtub3duQkVGTkhDK0FyaWFsLEJvbGRCRUZOSEMrQXJpYWwsQm9sZFZlcnNpb24gMC4xMUJFRk5IQytBcmlhbCxCb2xkVW5rbm93blVua25vd25Vbmtub3duAE8AcgBpAGcAaQBuAGEAbAAgAGwAaQBjAGUAbgBjAGUAQgBFAEYATgBIAEMAKwBBAHIAaQBhAGwALABCAG8AbABkAFIAZQBnAHUAbABhAHIAQgBFAEYATgBIAEMAKwBBAHIAaQBhAGwALABCAG8AbABkAEIARQBGAE4ASABDACsAQQByAGkAYQBsACwAQgBvAGwAZABWAGUAcgBzAGkAbwBuACAAMAAuADEAMQBCAEUARgBOAEgAQwArAEEAcgBpAGEAbAAsAEIAbwBsAGQAVQBuAGsAbgBvAHcAbgBVAG4AawBuAG8AdwBuAFUAbgBrAG4AbwB3AG4AAAADAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAsVSAQQ0DrACvA6wAAgAQA6wAIAOsAKADrAADAEADrLMHDTJAuAOssxIUMkC4A6yyFisyuf/AA6yyOjNAuAOssy2UMoC8A6sAXwAz/8ADq7JVM0C4A6uzQEQyQLgDq7MzOzJAuAOrsy8xMkC4A6uyCDNAuAOrswcUMh9BGgOrAC8DqwACAA8DqwAvA6sATwOrAI8DqwCfA6sAvwOrAAYAEAOrAN8DqwD/A6sAAwOoA6KyRh9AuAOlsggzD0EUA6UAAQBAA6UAzwOlAP8DpQADACADpQCvA6UA7wOlAP8DpQAE/8ADo7MJDDJAuAOjsggzD0EbA6MAAQAPA6MAEAOjAIADowCvA6MAzwOjAAUAbwOjAJ8DowD/A6MAAwCfA6IArwOiAAIDogOhshAfEEEKA54AfwOeAAIDmgAPAQEAH//AA5izEBQyQLgDmbMPEzJAQRADlQBQA5UAAgCwA00AwANNAAIAbwORAH8DkQAC/8ADS7ItMTK5/8ADS7MKDjIQQRADiwAgA4sAgAOLAAMAoAOLAAEAIAOLAEADiwAC/8ADi7MTFjJAuAODsg8RMrn/wAN7sjA0Mrn/wAN7sxAYMlBBFAN4AAEDZQNuACMAHwN+A24AHgAfA2MDbgAdAB8DYgNkAA0AH//AA0CzDxAygEEQAz8AAQM/AxUAKQAfA0EDFgAyAB8DRAMaABsAH//AA3WyDhEyuf/AA3WyKCoyQQoDQwMYADIAHwMPAw0ANAAfAwgDB7IyHyC7A0AAAQBAA4izCQsyQLgDiLIQFTK9A4UDBwAUAB8DgAMHshcfD70DCgAvAwoAAv/AA1SzCQ0ykEEMA1QAoANUAAIAHwNuAAEAnwNuAAEAQANusgkLMkERA0UDHAAWAB8DawMdABUAHwNGAx4AFQAfA6cDoQBGAB8DnbMmHB/AuwOTAAEAQAOSswkNMkC4Az6yCDNAuAM+sw0OMsBBCQM+AAEAsAOOAMADjgAC/8ADkLMmODIAQSYDKAAwAygAAgAgA38AMAN/AAIAEAOKADADigBQA4oAbwOKAH8DigCfA4oABgAAA4kAMAOJAAIALwN6AHADdwCQA3cAnwN6AAT/wAMVsg8QMrn/wAMVsiQoMrkDGQMYsjIfELsDGgAB/8ADGrMJDjJAuAMYshITMrn/wAMYswwOMj+9A3MATwNzAAIAQAN0sxcYMm+7AyoAAQBAAyyzGBsyQLgDcLIJDDK9AxcDFgAyAB//wAMWsg4RMr0DHAMeABYAHwMdAx6yFR+wQR8DHgABAA8DHwABAsoC0AAVAB8C0wLVAA0AHwLPAtAADQAfAssC0AANAB8CzQLQAA0AHwLOAtAADQAf/8AC0LMJDDJAuALSswkMMuBBHALlAAEAXwLdAJ8C5QACArsCwwAwAB8C2gK4ADIAHwLZArkAPwAfAtgCuABkAB8CuQK4ADMAHwK6siHIH7gCuLMhyB9AuAObsg0WMrn/wALDsisvMrn/wALDsh8lMrn/wALDshcbMrn/wALDshIWMkElAsICwQAcAB8C1wLBACQAHwLBAsAAIgAfAr8CwAAYAB8CwAJ0AMgAHwK1AjUAOwAfArQCNQA7AB8CxAK8AB4AHwK3ArYAOAAfArOyDsgfuAKwsgfIH7gCr7IGyB+4Aq6yAMgfuAKvslAvH7wCrgKrABoAHwKtsiYaH7gCqLMmJB8PuwI1AAECpQJ0sh0fEkEKAqEBWAH0AB8CoADYAfQAHwASAqKyN8gfuAKQsrwgH7kCkAKQQBg3QCVALUCmAzAlMC0wpgMgJSAtIDcgpiBBEAKOAAUAnwKLAAECiwKLADcAIAKJADACiQBAAokAkAKJsgQ3sEH9AnQAwAJ0AAIAgAJ0AKACdAACAGACdABwAnQAAgAAAnQAEAJ0AAIAgAJ0APACdAACAD8ChQBPAoUAAgCQAn4AkAJ/AJACgACQAoEABACQAnoAkAJ7AJACfACQAn0ABACQAnQAkAJ1AJACdwADAHACfgBwAn8AcAKAAHACgQAEAHACegBwAnsAcAJ8AHACfQAEAHACdABwAnUAcAJ3AAMAYAJ+AGACfwBgAoAAYAKBAAQAYAJ6AGACewBgAnwAYAJ9AAQAYAJ0AGACdQBgAncAAwBQAn4AUAJ/AFACgABQAoEABABQAnoAUAJ7AFACfABQAn0ABABQAnQAUAJ1AFACdwADAEACfgBAAn8AQAKAAEACgQAEAEACegBAAnsAQAJ8AEACfQAEAEACdABAAnUAQAJ3AAMAMAJ+ADACfwAwAoAAMAKBAAQAMAJ6ADACewAwAnwAMAJ9AAQAMAJ0ADACdQAwAncAAwAgAn4AIAJ/ACACgAAgAoEABAAgAnoAIAJ7ACACfAAgAn0ABAAgAnQAIAJ1ACACdwADABACfgAQAn8AEAKAABACgQAEABACegAQAnsAEAJ8ABACfQAEABACdAAQAnUAEAJ3AAMA4AJ+AOACfwDgAoAA4AKBAAQA4AJ6AOACewDgAnwA4AJ9AAQA4AJ0AOACdQDgAnexA9BBxQJ+ANACfwDQAoAA0AKBAAQA0AJ6ANACewDQAnwA0AJ9AAQA0AJ0ANACdQDQAncAAwAwAnQAQAJ0AAIAwAJ+AMACfwDAAoAAwAKBAAQAwAJ6AMACewDAAnwAwAJ9AAQAwAJ0AMACdQDAAncAAwCwAn4AsAJ/ALACgACwAoEABACwAnoAsAJ7ALACfACwAn0ABACwAnQAsAJ1ALACdwADAKACfgCgAn8AoAKAAKACgQAEAKACegCgAnsAoAJ8AKACfQAEAKACdACgAnUAoAJ3AAMAkAJ+AJACfwCQAoAAkAKBAAQAkAJ6AJACewCQAnwAkAJ9AAQAkAJ0AJACdQCQAncAAwAgAn4AIAJ/ACACgAAgAoEABAAgAnoAIAJ7ACACfAAgAn0ABAAgAnQAIAJ1ACACdwADAoEBWAgBAB8CgAEpCAEAHwJ/AOwIAQAfAn4A2AgBAB8CfQCxCAEAHwJ8AKYIAQAfAnsAgggBAB8CegA3CAEAHwJ3ACYIAQAfAnUAIAgBAB8CdAAfCAGyHzcPQRYCNQBPAjUAXwI1AG8CNQCfAjUArwI1AL8CNQAHAK8CNQDPAjUA3wI1AP8CNUAiBA8HTwefB68HvwcFrwfgBwIPBk8GnwavBr8GBa8G4AYCIEEbAg0AAQBfAjUAAQCPAjUAAQB/AjUA7wI1AAIALwI1AD8CNQACAD8CNABPAjQAAgI1AjUCNAI0QBHtIO8qAc8qAb8qAa8qAY8qAUEJAkcBBAAeAB8CIAA3AgEAHwFYQAwmPh/YJj4fNyYnPh+4Ao627BcfsiY2H7gBvLImNh+4ASlAKyY2H+wmNh+xJjYfpiY2H4ImNh83JjYfMiY2Hy0mNh8lJjYfHyY2HzcmKh+4AVhAIiY+H9gmPh+8Jj4fJyY+HyEmPh8gJj4fNwAWFgAAABIRCEC5Ag0BprPFDQAJuAG8sicoH7gBu7InMB+4AbiyJ08fuAG3sidiH0EJAbYAJwEBAB8BtQAgAqsAHwGvsh/kH7gBrbIf5B+4AayyH7sfuAGosh80H7gBXbInLh+4AVuyJ80fQQ0BVQAfBAEAHwFUAB8EAQAfAVMAHwIBAB8BUrIfVh+4AVGyHykfuAErsicmH0ENASoAJwElAB8BKQFYAOQAHwElAB8EAQAfASSyH+QfuAEjsh87H7gBIrIfOR9BDQEIACcIAQAfAQYALQEBAB8BBQAfAQEAHwEDsx+7H++5AVgEAUALH+0fkx/sH+Qf6x+4AgGyH9kguAQBsh/PJbgBVkAKH7wtnh+7H0EfskEKAVgEAQAfALEBWAQBAB8AsAFYBAG1H6YliR+buQFYASW2H5kfLh+OLbgIAbUfjR8pH4m5AVgEAbIfgiC4AqtAEx+AHzAfdC3kH3MfSh9hH1IfXSW4AquyH1wfvAgBAB8AWQFYAqu2H1AliR9JH7gBJbIfRyW4BAFACx9GH3kfQB8nHzkgvAKrAB8AOAFYBAGyHzctvAElAB8AMgFYASW2HywfNB8qJbgIAbIfVTe4ARFAKgfwB5AHWwdCBzsHIwciBx4HHQcUCBIIEAgOCAwICggICAYIBAgCCAAIFLj/4EArAAABABQGEAAAAQAGBAAAAQAEEAAAAQAQAgAAAQACAAAAAQAAAgEIAgBKALATA0sCS1NCAUuwwGMAS2IgsPZTI7gBClFasAUjQgGwEksAS1RCsDgrS7gH/1KwNytLsAdQW1ixAQGOWbA4K7ACiLgBAFRYuAH/sQEBjoUbsBJDWLEBAIWNG7kAAQEZhY1ZWQAYFnY/GD8SPhE5RkQ+ETlGRD4ROUZEPhE5RkQ+ETlGYEQ+ETlGYEQrKysrKysrKysrKxgrKysrKysrKysrGCsdsJZLU1iwqh1ZsDJLU1iw/x1ZS7CBUyBcWLkCDwINRUS5Ag4CDUVEWVi5BHACD0VSWLkCDwRwRFlZS7DkUyBcWLkAIAIORUS5ACcCDkVEWVi5CEIAIEVSWLkAIAhCRFlZS7gBJVMgXFi5ACYCD0VEuQAhAg9FRFlYuQoNACZFUli5ACYKDURZWUu4BAFTIFxYsdggRUSxICBFRFlYuSUAANhFUli5ANglAERZWUu4BAFTIFxYuQFYACZFRLEmJkVEWVi5IyABWEVSWLkBWCMgRFlZS7ApUyBcWLEfH0VEsS0fRURZWLkBDQAfRVJYuQAfAQ1EWVlLsC9TIFxYsR8fRUSxJR9FRFlYuQE1AB9FUli5AB8BNURZWUu4AwFTIFxYsR8fRUSxHx9FRFlYuRQoAB9FUli5AB8UKERZWSsrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKytlQisBszF1fsNFZSNFYCNFZWAjRWCwi3ZoGLCAYiAgsX51RWUjRSCwAyZgYmNoILADJmFlsHUjZUSwfiNEILExw0VlI0UgsAMmYGJjaCCwAyZhZbDDI2VEsDEjRLEAw0VUWLHDQGVEsjFAMUUjYURZsz88WEFFZSNFYCNFZWAjRWCwiXZoGLCAYiAgsVg8RWUjRSCwAyZgYmNoILADJmFlsDwjZUSwWCNEILE/QUVlI0UgsAMmYGJjaCCwAyZhZbBBI2VEsD8jRLEAQUVUWLFBQGVEsj9AP0UjYURZRWlTQgFLUFixCABCWUNcWLEIAEJZswILChJDWGAbIVlCFhBwPrASQ1i5OyEYfhu6BAABqAALK1mwDCNCsA0jQrASQ1i5LUEtQRu6BAAEAAALK1mwDiNCsA8jQrASQ1i5GH47IRu6AagEAAALK1mwECNCsBEjQgArKysrKysrKwCwEkNYS7A1UUuwIVNaWLEmJkWwQGFEWVkrKysrKysrKysrKysrKysrKysrc3Nzc3NFsEBhRBgARWlERWlEc3NzdHNzc3RzdHN0KysrKysrKysrKysrAHNzc3Nzc3Nzc3Nzc3Nzc3Nzc3Nzc3N0dHR0dHR0dHR0dHR0dHR0dHR0dHR1dXVzdHV1dXUrcwAAS7AqU0uwNlFaWLEHB0WwQGBEWQBLsC5TS7A2UVpYsQMDRbBAYESxCQlFuP/AYERZK0VpRAF0AHNzcytFaUQrAStDXFhACgAGAAcCoAagBwK5/8ACdLMaHTJvvQJ3AH8CdwAC/8ACd7IvMTK5/8ACd7MiJTJAuAJ0sy81MkC4AnSzKCoyQLgCdLIaITK4/8CzNxodMrj/wLMlGh0yuP/AQBEtGh0ykCWQLZA3oCWgLaA3Brj/wLamGh0yH6YfuAKOsi+mAwB0K3MrKysrKysrK3Qrc3RZACsrQ1xYuf/AAqGyHB0yuf/AAqCyHB0yKytZK3MBKysrKwArKysrKysrKysrKysrKysrKysBKysrKysrK3N0KysrKysrKytzcysrKysrK3MrcysrK3QrKytzc3NzcytzcysrK3MrKwArKysrc3RzK3MrKysrdSsrKysrKysrdSsrKysrcysrKytzdHUrK3NzcysrK3Mrc3N0dSsrc3R1KytzdHUrKysrKysrKysrKyt0dSsAAA==); }&#xA;@font-face { font-family: &quot;g_font_2&quot;; src: url(data:font/opentype;base64,AAEAAAANAIAAAwBQT1MvMmJoWKEAAADcAAAATmNtYXCjekLVAAABLAAAAIhjdnQgoRzX6wAAAbQAAAZUZnBnbcx5WZoAAAgIAAAGbmdseWb07S6AAAAOeAAAcspoZWFk5t1y1gAAgUQAAAA2aGhlYRIzFiYAAIF8AAAAJGhtdHh0wP1UAACBoAAANXRsb2NhBeMkhgAAtxQAADV4bWF4cBK5AcEAAOyMAAAAIG5hbWU0cTvsAADsrAAAAi5wb3N0AAMAAAAA7twAAAAgcHJlcCXWTb8AAO78AAALvgAABAABkAAFAAAEAAQAAAAEAAQABAAAAAQAAGYCEgAAAQEBAQEBAQEBAQAAAAAAAAAAAAAAAAAAAAA/Pz8/AEAAIACpCAACAADMCAwDmAAAAAAAAQADAAEAAAAMAAQAfAAAABoAEAADAAoAIAAlACkAOgA9AD8AWQBfAHoAqSAZ4AH//wAAACAAJQAoACsAPQA/AEEAXwBhAKkgGeAA////4//j/+P/4//j/+P/4//j/+P/4uCdAAAAAQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAABAAAAAMAEAW6ABkFugAaBacAGQQmABgAAP/nAAD/6AAA/+f+af/oBboAGf5p/+gC6gAAALgAAAC4AAAAAACoAK0BaQCtAL8AwgHwABgArwC5ALQAyAAXAEQAnAB8AJQAhwAGAFoAyACJAFIAUgAFAEQAlAEZ/7QALwChAAMAoQDNABcAVwB+ALoAFgEY/+kAfwCFA9MAhwCFAA0AIgBBAFAAbwCNAUz/dQBcAN8EgwA3AEwAbgBwAYD/WP+O/5L/pAClALkDyP/9AAsAGgBjAGMAzf/uBdj/3AAtAFwAlQCZAN8Bkgm1AEAAVwCAALkDnQByAJoDXQQB/2f/+gADACEAdwDNAAQATQDNAcACKwBMAGUA5wEYAXwDQwXY/6P/sP/EAAMAHABdAGgAmgC6ATUBRwIhBVz/Tf/NABYALQB4AIAAmQCyALYAtgC4AL0A2gEMBfD/pP/wABkALABJAH8AtADOAcAD/v2B/j8AAAAFABgAKQA5AEkAbwC+AMcA0AEjAcECbwUMBTIFQAV6/9QAFAAxAFUAVwCnALQA5gH3An4CfgJ/A8YERv9CAA4AhQCRAL8AwgDFAOEBGgEvAU8BVgIpAm8CngNyAAgALAAxADEAZABpAIkAmADHAN4BKwG2AgwCzwOjBKsE+wYd/uD/DgAGACYAmwCdAMEBDQEYASABcwGCAdYB4wJDAl8CmwLiA5QEqQTSB2EAHABeAG0AjQCrAPcBEgE4AVEBWwFoAXwBhwGRAZkBzQHQAegCQQJUAmsC7wNoA3EDvQRCBEIEUwRzBIMFhgWLBuj+WP7E/tH+9/8y/4YAUQB8AIEAkQCVAJ4AtAC5AM8A2QDZAN8A4gEFAQsBDgEOASABIQFVAXsBewF+AY0BogGoAakBtAHQAdAB4gHpAfIB9QH7AgACAAIGAhsCIQIiAiICIwJyAncClAKcAs8CzwLQAuwC+QMXAyIDKwM1AzwDWQNvA3EDhwOQA5ADtQPhBBoEzwT/BTIFMgWWBZ8FqAWrBcIF8AYMB4IIAAjM/KP9Kv3e/gD+iP6W/rL+tP/hABUAGQAaABwAHwA8AFEAYQBhAGoAeACWAKUArwDTAQwBGAEaASoBPgFMAVEBXwFqAXEBeAGCAYQBmgGlAagBqQGuAbwBzQHXAe8CAAINAhwCIQIiAi4CNQJCAk8CTwJeAmUCcQKQApICtALWAvoDBwMLAw8DFQMqA0cDXQNlA3QDeQOWA7ADzAPdA+ID9gP8A/wD/wQKBB8EIgQmBCsERwRfBHUEngTnBOcFXAXLBeUGCgZtBoYGuAbxBzYHPgdQB1EHXQePB7YH1AhgALYAwwC1ALcAAAAAAAAAAAAAAAAB4AOBA0UDtQCOAjMEGQLOAs4ALQBfAGQDTQI/AAACqAGIAn0BtAIkBXgGOwI7AU4A8AQmApQCxgKfAvYCOwNNAUsBUwBqAjEAAAAAAAAGFASqAAAAPATDAO0EvAJlAs4DtQB4BgwBfgLvBgwAsgEAAjkAAAHFAzAEKwPLANoD3wEHBKEA2wQKARcB7QKnA1ABCwG9BD4FWAAhA5wArgNxAX0AtQJFAAAK+wiMASsBTgGqAIcAVAEyAfgD/wADAk4AtAA3A+MAgwBrAtgA7QB3AIgAlwFkBGcAjgAzAXwA5wCmAp4DKQVuBioGFQHJAmkEigITAbQAAgSpAAACOQEkAQMFFACEAV0DmgbvAtkAdQDPBAoA3gOsBLwCzwKuA00E8AVSAWgAbQB9AIYAcf+BAHkFWATSAWcAAwFWACUE4ACUAHwDMgQhAJQAfwByAFwALwC2ABgAugC4AEEDTQByABgAHwBMAWoBVQCZAJoAmgCYALIABAB4AGkAFABXAG4AzgC0BlQCuABnBQ4BZQDnAAAEy/5SAFr/pgCZ/2cAbv+SAC3/1ACH/3wAuACoAOUAjwCoAYX+ewBwAB4A2QDeAUwFRgLPBUb/LQKKAtkCUwKWALcAAAAAAAAAAAAAAAAAAAElARgA6gDqAK4AAAA+BbsAigTXAFMAP/+M/9UAFQAoACIAmQBiAEoA5ABtAO4A5QBIA8AAM/5OArH/RgNwAHkF3wBR/6f/HwEKAGj/bABPALwApQcFAGEHKwDtBLAB0gC2AHsAZQJS/3QDZf5pAJQAjwBcAEAAhgB1AIkAiUBDVVRBQD8+PTw7Ojk4NzU0MzIxMC8uLSwrKikoJyYlJCMiISAfHh0cGxoZGBcWFRQTEhEQDw4NDAsKCQgHBgUEAwIBACxFI0ZgILAmYLAEJiNISC0sRSNGI2EgsCZhsAQmI0hILSxFI0ZgsCBhILBGYLAEJiNISC0sRSNGI2GwIGAgsCZhsCBhsAQmI0hILSxFI0ZgsEBhILBmYLAEJiNISC0sRSNGI2GwQGAgsCZhsEBhsAQmI0hILSwBECA8ADwtLCBFIyCwzUQjILgBWlFYIyCwjUQjWSCw7VFYIyCwTUQjWSCwkFFYIyCwDUQjWSEhLSwgIEUYaEQgsAFgIEWwRnZoikVgRC0sAbELCkMjQ2UKLSwAsQoLQyNDCy0sALAXI3CxARc+AbAXI3CxAhdFOrECAAgNLSxFsBojREWwGSNELSwgRbADJUVhZLBQUVhFRBshIVktLLABQ2MjYrAAI0KwDystLCBFsABDYEQtLAGwBkOwB0NlCi0sIGmwQGGwAIsgsSzAioy4EABiYCsMZCNkYVxYsANhWS0sRbARK7AXI0SwF3rkGC0sRbARK7AXI0QtLLASQ1iHRbARK7AXI0SwF3rkGwOKRRhpILAXI0SKiocgsKBRWLARK7AXI0SwF3rkGyGwF3rkWVkYLSwtLLACJUZgikawQGGMSC0sS1MgXFiwAoVZWLABhVktLCCwAyVFsBkjREWwGiNERWUjRSCwAyVgaiCwCSNCI2iKamBhILAairAAUnkhshoaQLn/4AAaRSCKVFgjIbA/GyNZYUQcsRQAilJ5sxlAIBlFIIpUWCMhsD8bI1lhRC0ssRARQyNDCy0ssQ4PQyNDCy0ssQwNQyNDCy0ssQwNQyNDZQstLLEOD0MjQ2ULLSyxEBFDI0NlCy0sS1JYRUQbISFZLSwBILADJSNJsEBgsCBjILAAUlgjsAIlOCOwAiVlOACKYzgbISEhISFZAS0sS7BkUVhFabAJQ2CKEDobISEhWS0sAbAFJRAjIIr1ALABYCPt7C0sAbAFJRAjIIr1ALABYSPt7C0sAbAGJRD1AO3sLSwgsAFgARAgPAA8LSwgsAFhARAgPAA8LSywKyuwKiotLACwB0OwBkMLLSw+sCoqLSw1LSx2uAIjI3AQILgCI0UgsABQWLABYVk6LxgtLCEhDGQjZIu4QABiLSwhsIBRWAxkI2SLuCAAYhuyAEAvK1mwAmAtLCGwwFFYDGQjZIu4FVViG7IAgC8rWbACYC0sDGQjZIu4QABiYCMhLSy0AAEAAAAVsAgmsAgmsAgmsAgmDxAWE0VoOrABFi0stAABAAAAFbAIJrAIJrAIJrAIJg8QFhNFaGU6sAEWLSxLUyNLUVpYIEWKYEQbISFZLSxLVFggRYpgRBshIVktLEtTI0tRWlg4GyEhWS0sS1RYOBshIVktLLATQ1gDGwJZLSywE0NYAhsDWS0sS1SwEkNcWlg4GyEhWS0ssBJDXFgMsAQlsAQlBgxkI2RhZLgHCFFYsAQlsAQlASBGsBBgSCBGsBBgSFkKISEbISFZLSywEkNcWAywBCWwBCUGDGQjZGFkuAcIUViwBCWwBCUBIEa4//BgSCBGuP/wYEhZCiEhGyEhWS0sS1MjS1FaWLA6KxshIVktLEtTI0tRWliwOysbISFZLSxLUyNLUVqwEkNcWlg4GyEhWS0sDIoDS1SwBCYCS1RaiooKsBJDXFpYOBshIVktLEtSWLAEJbAEJUmwBCWwBCVJYSCwAFRYISBDsABVWLADJbADJbj/wDi4/8A4WRuwQFRYIEOwAFRYsAIluP/AOFkbIEOwAFRYsAMlsAMluP/AOLj/wDgbsAMluP/AOFlZWVkhISEhLSxGI0ZgiopGIyBGimCKYbj/gGIjIBAjirkCwgLCinBFYCCwAFBYsAFhuP+6ixuwRoxZsBBgaAE6LSyxAgBCsSMBiFGxQAGIU1pYuRAAACCIVFiyAgECQ2BCWbEkAYhRWLkgAABAiFRYsgICAkNgQrEkAYhUWLICIAJDYEIASwFLUliyAggCQ2BCWRu5QAAAgIhUWLICBAJDYEJZuUAAAIBjuAEAiFRYsgIIAkNgQlm5QAABAGO4AgCIVFiyAhACQ2BCWblAAAIAY7gEAIhUWLICQAJDYEJZWVlZWS0ssAJDVFhLUyNLUVpYOBshIVkbISEhIVktAAAAAgEAAAAFAAUAAAMABwAAIREhESUhESEBAAQA/CADwPxABQD7ACAEwAAABQB3/8oGnwXTAAsAFwAbACcAMwEHQAqQGZAaAmgIGhsbuAKaQA8YGRQYGBkYGxUPGRoxKxK8Ap8ACQFlAAwCn0ALAxoZGQMBGxgYJSi8Ap8AHwFlAC4Cn7IlCxy8ApoAKwEAADECmrMirDUGvAKaABUBAAAPAppACSAAAQB1NFdaGCsQ9l3t9O0Q9u307QA/7f3tEDwQPD88EDwQ7f3tARESOTkREjk5hy4rfRDEMTAYQ3lAUgEzKR4rHwAzIDEfAS0mKx8ALyQxHwENAg8fABcEFR8BEQoPHwATCBUfASodKB8BMiEoHwEsJy4fADAjLh8ADgEMHwEWBQwfARALEh8AFAcSHwAAKysrKysrKysBKysrKysrKyuBAV0TNDYzMhYVFAYjIiYBIgYVFBYzMjY1NCYDATMBATQ2MzIWFRQGIyImASIGFRQWMzI2NTQmd56WirW3hoWxATlDWVpCRFlaQgMikvzhAeWel4q1t4eFsQE6RFlaQkVZWgRandzFv7rJxgHFdJuNc3SajnP6cwYJ+fcBjp7bxb+6yccBxHSbjHR0mo5zAAEAfP5RAmAF0wAQAD1ACicPAQAQEgcIEBC4ATOzAJ8OCLgBM0ARB58OXgADEAMgAwMDrBGdjBgrEPZd/fbtEPbtAD88PzwxMAFdASYCETQ3NjczBgcGBwYVEAEB35XOTVq8gXknPSMrASv+UbwB+AEO7tr9+9BZipa7vf4f/iAAAQB8/lECYAXTABAAZUAMKAIoEAIJChABABIJuAEzswqfAwG4ATO0AJ8DXg64//C0EBACVQ64//i0Dw8CVQ64/+S0DQ0CVQ64/+xADwoKAlUPDh8OAg6sEp2MGCsQ9l0rKysr/fbtEPbtAD88PzwxMAFdEyMAETQnJicmJzMWFxYVEAL9gQErKyI9J3qBvFpNz/5RAeAB4by5lopa0vv92u7+8v4IAAEAcgDtBDoEtgALADhAHwBuCQL5CANuBQcGCW4KBAr5BQFuPwJPAgICGQxXWhgrThD0XU30PO08EOQ8PAAv9Dz9PPQxMCURITUhETMRIRUhEQIB/nEBj6oBj/5x7QGSqAGP/nGo/m4AAQCq/t4BgwDNAAoATrUKAwAHqwa4AVBAJgEDPAICAQoBPAAKAgMBAzwABjgHOk8AXwBvAH8AoAAFAKALoZgYKxD0XfTkEO08EDwAP+08EDwQ7RD97QEREjkxMDM1MxUUBgcnNjY3ts1QVzI5NgPNzXGLJk0ZYVsAAQBBAbgCagJtAAMALEAZcAJwAwJNAU0CAgEjAAIaBXAAAQAZBHCNGCtOEORdEOYAL03tMTAAcQFdEzUhFUECKQG4tbUAAAEAugAAAYcAzQADACVAGAI8AAoCPF8AbwB/AK8ABKAAAQCgBKGYGCsQ9l1d7QA/7TEwMzUzFbrNzc0AAAEAAP/nAjkF0wADAFO5AAP/3rIUOQK4/95AIBQ5lwMBAgOfA68DAgN2AAEUAAABAgEAAwAKA+gAAugBuAGptQAABLN6GCsQPBD07RDtAD88PzyHBS4rXX0QxDEwAV0rKxUBMwEBqZD+WBkF7PoUAAACAFX/5wQRBcAAEAAdAVWxAgJDVFhAChoeBAUUHg0NFwm4/+i0Dw8CVQm4/+hAGQ0NAlUJEQAMDw8CVQAWDAwCVQAMDQ0CVQAvKysrzS8rK80AP+0/7TEwG7EGAkNUWEAKGh4EBRQeDQ0XCbj/9LQPDwZVCbj/5rQNDQZVCbj/7kAZCwsGVQkRABANDQZVABAMDAZVABALCwZVAC8rKyvNLysrK80AP+0/7TEwG7QGIBkQHLj/8LICIAu+/+AAFv/gABL/4AAP/+BAYgQGhwKIC4gPyQ4FCQcLGAJFE0wVShlDG1QTXBVcGVIbawdrC2MTbBVrGWAbeQJ3BnYLeg+HBpgHlhDJGNoC1gbWC9sPGhoeBAUUHg0NF3MJQCEjNDAJAQAJEAkCCZAfEXMAuP/AQA4hIzQgAEAAAgCQHseLGCsQ9l0r7RD2XXEr7QA/7T/tMTABXXEAXQA4ODg4OAE4ODhZWRMQEjYzMhYWEhUQAgYjIicmExAWMzI2ERAmIyIHBlVr06B2snRCatOh1HmRual8fKmpfnxKXQLTAQQBPaxfs/7/2v7+/sOtmLcBnf6X7/ABaAFq7mmGAAABAN8AAAL7BcAACgCvQCADQA0RNGsEfwKPApkIBKwEAQkABgUCAwkFAQwCAcoKALj/wEAKISM0MAABIAABALj/4LQQEAJVALj/6kARDw8CVQAcDAwCVQAODQ0CVQC4//BAGQ8PBlUAEAwMBlUAEA0NBlUAGgwFQA0PNAW4/8BADiEjNDAFASAFQAUCBRkLugE8AYUAGCtOEORdcSsrEPYrKysrKysrXXErPE39PAA/Pxc5ARE5MTABXQBdKyEjEQYGBzU2NjczAvu0QdNUl+IvdAR7PnwfrkfKXwAAAQA8AAAEBwXAAB4Bx7EGAkNUWEAJERANGBMTBlUNuP/0tBERBlUNuP/uQAkQEAZVDR4UBR64/+hAFxMTBlUeHhERBlUeHA4QBlUeDA0NBlUeuAK7QAwCChcXIB8QEQICIB8REjkv1M0REjkvzQAv7SsrKys/7SsrK8QyMTAbsQICQ1RYQAkREA0MEhICVQ24//RACQ8RAlUNHhQFHrj/4EALEhMCVR4UDxECVR64AruyAgoXuP/otAsLAlUXuP/sQA4NDQJVFxcgHxARAgIgHxESOS/UzRESOS8rK80AL+0rKz/tKyvEMjEwG0A2OwU7BrsFvwa7B8cIyRwHSQxZDFQOawxkDnoSehOJErwS5RrlG/AaDL8LtxMCGxAcEB0QHhAGvv/wAAf/4AAI//AACf/wQBoeChAIBgbKHBoUHBwaCBwaAwECCBocAw0eELgCpLNPEQERuAEYtQ0eFAUAHrgCu0APAQIMCnMX0wAAAUAhIzQBuwKBACAAEAE4QAwRtT8CXwJvAn8CBAK6AiQAHwGPsYsYKxD2XfTtEPYrPBD07QA/PP08P+39XeQREhc5ARESFzmHDi4rDn0QxAEREjkxMAA4ODg4ATg4ODgAXQFdcllZJRUhJjc2Njc2NjU0JiMiBgcnNjYzMhYVFAYGBwYGBwQH/DcCFyWjmu+omXuCnAG5E/jR0/ZIp8KiXB6trUE8Y8B+xOVma5OcihPP2eqtWKq8pIhhMQABAFb/5gQWBcAAKwFZsQICQ1RYQAsZGEANDQJVGBwAAbj/wEArDA0CVQEpIwoNDwwPHgoKKRUeHAQeKRwFKQ0jDQwYGQEAEiAQDAwCVSAHJrj/6LQMDQJVJi8rzS8rzS/NL80vABI5Pz8Q7RDtEjkv7cYQxhI5EMQrMhDEKzIxMBtAKAUNFg1FDYYNBEURVxF2GwNSFmwQahRkFnUNeRSGDYoUiRulDQoFIAO4/+BACwsMDQ4EBwEjDQwBuAKks0AAAQC7ARgAKQANATW0DAwVBBi6AqQAGQJoQCcVHhwFBB4pDRJzXyBvIAIgGA0NBlUggAdzJkAhIzQwJgEAJhAmAia4//S3DQ0GVSaQLRi4ATiyGdMBugE4AAD/wEALISM0IABAAAIAkCy4AZKxixgrEPZdK+307RD2K11xK+30K13tAD/tP+395BESOS/tEP1d5BESOQEREhc5MTABODgBXQBdAXFZEzcWFjMyNjU0JiMiBzcWMzI2NTQmIyIGByc2NjMyFhYVFAYHFhYVFAAjIiZWtB+Va3+von0zTBQSC3O4hmppjBS0IequeMprZmSCkP7o1sH/AYMYmYewgnyhFJ4CeH1jgoSEILXHZ7JkX5wuHr2OwP715gACABoAAAQQBboACgANASZANhJYDGgMmgypDMkMBUwDTA2UBAMSAQIIAAwGAwcFCgsDBwAMDA0NygMEFAMDBAMNAAIMDQQHA7sCuwAIAAIBoEAKAAQEAAwMAMoKBLgCZrcFBQpAHR80Crj/4LQQEAJVCrj/5rQNDQJVCrj/7rQNDQZVCrgBN0ANB0AiIzQHgCE1B5APArj/wEALDRQ0AAIQAiACAwK4/+C0DQ0CVQK4/+S2DQ0GVQK1DrgBjLGLGCsQ7CsrXSsQ9isr9CsrKys8EOYQ/TwAPz8Q9Dz2PBE5OQEREjk5hy4rBH0QxA8PDzEwAUNcWLkADf/eshI5Dbj/1EALMzkDIi05AwQdHTwrKysrWV0AXUNcWEAUDEALOQyAUDkMQCY5DCIcOQxALTkrKysrK1khESE1ATMRMxUjEQMRAQKW/YQCnZPGxrT+NQFfpQO2/Eql/qECBAKV/WsAAQBV/+cEIQWmAB4BVrECAkNUWLkAAf/AQA0NDQJVARwOCh4VFRwSuAK7QAsPBAQeHA0OAQAHGLj/6rQPDwJVGLj/6rQNDQJVGC8rK80vzS8AP+0/7RI5L/3EEMQrMTAbQCkSDA0NBlUPDA0NBlVLGnkdih2WE6cTwwzWDNsbCAkTGA4qGgMJMAUwC7r/4AAD/+BAEBMKFRITE8oODxQOExQODw24AqRAEw4KHhVADqAOAg4OD0AVARUVHBK4Aru3DwQB00AAAQC4ARhAIAQeHA0RXxBvEH8QjxAEEIAHcxhAISM0MBgBABgQGAIYuP/0tw0NBlUYkCASvAE1AA8BlQANATiyDrUBugE4AAD/wEALISM0IABAAAIAkB+4AZKxixgrEPZdK+307fTtEPYrXXEr7fRdPAA/7f1d5D/tEjkvXRE5L10Q7RDkhwguKwV9EMQAERI5MTABODg4OAFxXSsrWRM3FhYzMjY1NCYjIgYHJxMhFSEDNjMyABUUBwYjIiZVvRWZbIK0rYxXjCipjgLZ/bdPhJHAAQh0jfTI/QGAEIqLxKKask8/FgLxrP52XP720ceRsuAAAAIATf/nBBUFwAAdACoBT7ECAkNUWEAfDwEfAV8BAwEbKB5ADQENDRQFHhsFIh4UDQoeAQAlELj/9EAZDQ0CVRAeFxAPDwJVFxAMDAJVFwwNDQJVFy8rKyvNLyvN1M0QxQA/7T/tEjkvXe0QxF0xMBtALWsZAUQHQBVEGUQgWhJUIGsDZAdkCGoSZCB0CHUchQiGHNYI1BYRByANDQZVJ7j/4LQNDQZVI7j/4EALDQ0GVSEgDQ0GVQe4/+C0JyAjICG4/+BAESgeQA1QDQINDRQbAdNfAAEAuAJoQAkFHhsFIh4UDQG4AThAEgC1JXMQQCEjNDAQAQAQEBACELj/8LcMDAZVEJAsCroBOAAeATlAFj8XXxdvF38XBBcWDAwGVRcWDQ0GVRe4AiSzK8eLGCsQ9isrXe3tEPYrXXEr7fTtAD/tP+39XeQREjkvXe0xMAE4ODg4KysrKwFdAF1ZAQcmJyYjIgcGBgc2NjMyEhUUBgYjIgAREDc2MzIWARQWFjMyNjU0JiMiBgP7sxgsSWtWQVViAkG8Z7T9d9CE4f7knYnord39N0+OTnKkont6qgRTDmowTTA+7txjYP730ortfgFLAXwBqcGowvzdXapZuJ6Yr68AAQBhAAAEFgWnAA0AcEAOxA0BBA0BBAIIBAkDDQC4ArtAMAIBBAkMDXMDAwJAISM0TwJfAm8CAwIaDwhzCesATwFfAV8CAz8BXwFvAX8BBAEZDrgBkrGLGCtOEPRdcTxN9O1OEPZxKzxNEO0APz88/Tw5ETkBERI5MTABcV0TNSEVBgADBgcjNhISN2EDtYz+7Us2D7kDgvOJBPqtjJX+Ev77uNutAeoBx5wAAAMAU//nBBkFwAAXACMAMAIAsQICQ1RYtAwAGx4uuP/AQBcTEwJVLi4SIR4GBSgeEg0eCQwMDAJVCbj/9LYNDQJVCSsPuP/wtA8PAlUPuP/otAsLAlUPuP/otg0NAlUPGAO4//C0EBACVQO4//C0Dw8CVQO4//RAGQ0NAlUDJBUMCwsCVRUMDAwCVRUMDQ0CVRUvKysrzS8rKyvNLysrK80vKyvNAD/tP+0SOS8r7Tk5MTAbsQYCQ1RYtx4JDAwMBlUJuP/0tg0NBlUJKw+4/+S0Dw8GVQ+4/+S2DQ0GVQ8YA7j/8LQPDwZVA7j//EAiDQ0GVQMkFQwMDAZVFQwNDQZVFQwAGx4uLhIhHgYFKB4SDQA/7T/tEjkv7Tk5AS8rK80vKyvNLysrzS8rK80xMBtANzUWASkWSRZJJuYM6TAFCTABfQB9AXwEdAhxC3IMdQ16F4sAigGMBIYIgQuEDIYNjRfMEcYTEiK4/+CyHCAauP/gsiAgL7j/4LItICa4/+BAHikgDAAeGAAMGx4uoC4BLhIhHgYFKB4SDR5zvwkBCbgCZ0AQK3MPQCAjNDAPAQAPEA8CD7gBkbYyGHOwAwEDuAJnsiRzFbj/wEAOISM0IBVAFQIVkDHHixgrEPZdK+30Xe0Q9F1xK+30Xe0AP+0/7RI5XS/tOTkBERI5OTEwATg4ODg4ODg4AV1ycQBxWVkBJiY1NDYzMhYVFAYHFhYVFAAjIgA1NDYTFBYzMjY1NCYjIgYDFBYWMzI2NTQmIyIGAWpwbOa/wOprbYeN/vbZ2f72kWKGa2iFiWZniDpJkFOBqK2Cf6cDGymYaqDa36BmlyksxIi8/wABAcCPwQFUaISDX2OHhPz/TZBPpoCCqqgAAAIAVf/nBBkFwAAeACoBrrEGAkNUWLcLHxgBACURGLj/9rQPDwZVGLj/9LQNDQZVGLj/8EAoDAwGVRgRDA0NBlUREAwMBlURGBEsKwsoHg8OHw5PDgMODhQAUAEBAbj/wEANEBEGVQEEHhwNIh4UBQA/7T/txCtdMhI5L13tMgEREjk5LysrLysrKxDN1M0Q3cUxMBuxAgJDVFi3Cx8YAQAlERi4/+q0Dw8CVRi4/+pAKg0NAlUYEQwMDAJVERgRLCsLKB4PDh8OTw4DDg4UAFABAQEEHhwNIh4UBQA/7T/txF0yEjkvXe0yARESOTkvKy8rKxDN1M0Q3cUxMBtANDoaTBZAI1sWVyNmA2wWbRpnI3oafR6MGosemhapGrwa6hbmIPYgEz0WnhatFgM6KWQGAie6/+AAI//gQBghIAYgKB5PDl8OAg4OHCIeFAUB01AAAQC4Ami0BB4cDR+6ATkACwE4QBEYQCEjNDAYAQAYEBgCGJAsAbgBOLQAtSVzEbj/wEAOISM0IBFAEQIRkCvHixgrEPZdK+307RD2XXEr7e0AP+39XeQ/7RI5L13tMTABODg4OABdcQFdWVkTNxYWMzI+AjU0JwYGIyICNTQAMzIWEhEQAgYjIiYBNCYjIgYVFBYzMjZwrRZ8YVN9UDYBNrtttvwBB8aP7Xt68aKs2gLLpXR4sql8faEBUxB6bkx/2HAMGFZrAQjY3wEQmv7j/vL+5/6zrr8DNJu2xJyMr68AAAIAuQAAAYYEJgADAAcAOEAgBAUABgcJAgY8BAM8AQYECgI8LwA/AAIgAAEAoQihmBgrEPRdce0APz/tEO0BERI5ORI5OTEwEzUzFQM1MxW5zc3NA1nNzfynzc0AAgByAaEEOgQGAAMABwBHQCcFBgEEBwkAJQMBJQMCByUEBAYlMAIBnwLPAgICvwUAGgkBGQhXWhgrThDkEOYAL03tXXHtPBDtEDztEO0BETk5ETk5MTABITUhESE1IQQ6/DgDyPw4A8gDXqj9m6gAAAIAWgAABAwF0wAeACIAhEAvjBqLGwJ8GnwbAmIaZRsCawxhDgJaDFQOAjYORA4CGxkIBwQAECcREQANKRQBHgC4Aq9AIyEiITwfCh88IiIgPCEhHgBeHm4KXhdqJBBeIBEBEWojV1oYKxD2Xe0Q9u307RA8EO08EP0AP+08EPY8P+0SOS/kERc5MTABXV1dXQBdXQEmNTQ3Njc+AjU0JiMiBgcnNjYzMgQVFAYHDgIHAzUzFQHYAR4WMSS7OKR3c5oYuRn3y9cBAFqDWDYaArjNAWkkEmpNOjsrpWI6aZ+QmRbN2uqmYKJ0TkpgbP6Xzc0AAv/9AAAFWQW6AAcADgFntgEODxACVQK4//K0DxACVQK4//i0DQ0GVQK4//RAWQwMBlUJDAwMBlUFDAwMBlUvEDAQZwhoCWAQiAOQEMkFxgbAEPAQCwgFWQFWAlAQaAuwEPMM8w3zDgkEDAQNBA4DCwoJBQQEDA0OCAYHBwwJBQQIBgwHAQAAuP/4QA8MDAJVACAHDBQHBwwCAwO4//hAFQwMAlUDIAQMFAQEDAkeBQUIHgYDBrgCcEAJAAgM6UACAQICugELAAEBC0ASDCAAZQcDUlAEzwTfBAOQBAEEuAEBQAtQDMAH3wwDkAwBDLgBAUAQDwfPBwJ/B4AHAgeTD9bXGCsQ9F1xGfRdcfRdcRjtEO0aGRDt7QAYPzwa7T/kPBDtPBDthwUuKyt9EMSHLhgrK30QxAEREjk5ETk5hxDExA7ExIcFEMTEDsTEMTABS7ALU0uwHlFaWLQEDwMIB7r/8AAA//g4ODg4WQFycV0rKysrKysjATMBIwMhAxMhAyYnBgcDAjPRAljdq/2bodkB8ZlGIhwzBbr6RgG8/kQCWgGWuXeNiwAAAwCWAAAE6QW6ABEAHQAqARO5AAT/9EBHCwsGVQQERiNWI2YjcwmECQZpGnUFcAlzC4MFgwsGJxYJAxgnKh4WHQkJExIeKiopKQAcHR4CAQIfHh4RAAgYJgYMEBACVQa4/+ZAMw8PAlUGEg0NAlUGBgwMAlUGCAsLBlUGDAwMBlUGFA0NBlUGVCUmDBwQEAJVDAoNDQJVDLj/9EAVCwsGVQwaLB0eIAEgAAEAIBAQAlUAuP/2tA8PAlUAuP/2tA0NAlUAuP/6tAwMAlUAuP/6tAwMBlUAuP/wQAoNDQZVAF0rO1wYKxD2KysrKysrXTz9PE4Q9isrK03t9CsrKysrKyvtAD88/Tw/PP08EjkvPBD9PDkvETkREjkBEhc5MTABXQBdKzMRITIWFhUUBgcWFhUUDgIjASEyNzY2NTQmJiMhESEyNz4CNTQmJiMhlgImqMtzZmeFj1eAwYz+kwE9gThKS0aCnv7bAW1eJkNaOlSVjP6tBbpZuWVepjMnvIBnsWAxA1IRFmZNSW8p+6AHDDhrRlJ5MQAAAQBm/+cFdgXTAB0A07VjAmodAgG4/+i0CwsGVQC4/+hAXwsLBlUgADINYwBwAHQdgACEHZAAmgWrA6UNuQO0DccN0ADkHfMdEQ4SHREdHQMqBigRKhwgH0cNVhRXFVYZaAVrHXsSixKaA5kOmhyoAaQCqBHVDhMAFAAaEBQQGgQCuP/esig5Abj/wEAtKDkQDwABBBsTHgwDGx4ECRAmD0oAJiABAQEaHxcmIAgBCAwLCwZVCBkeY1wYK04Q9CtdTe1OEPZdTe307QA/7T/tERc5MTABKytdXXEAXSsrAXIBFwYEIyIkAjU0EiQzMgQXByYmIyIGAhUUEhYzMjYEtMI9/sPl7f7Xm68BQ8LcASw7vzPCk6njXG3mhqPiAgIx7/vBAW7S5QFVseDLLaCSov7vkbv+6Yq8AAACAJ4AAAVaBboADwAdAOVALyAfAUMIHB0eAgECERAeDwAIFyYgCQEfQA0NAlUJIBAQAlUJCg8PAlUJGA0NAlUJuP/0QBUMDAZVCRofHRAgASAAAQAgEBACVQC4//a0Dw8CVQC4//a0DQ0CVQC4//q0DAwCVQC4//e0DAwGVQC4//hACg0NBlUAXR47XBgrEPYrKysrKytdPP08EPYrKysrK13tAD88/Tw/PP08MTBDeUA2AxsHCAYIBQgECAQGGRgaGAIGCwoMCg0KAwYVFhQWExYDBhsDFyEBEg4XIQEYCBwhARYKESEAKysBKysqKioqgQFdMxEhMhcWFxYSFRQCDgIjJSEyNjc2NjU0JicmIyGeAfmrWn5ZdHNOepHNhf6xATmRpTFFTZdsTq3+zAW6FR1MYv7PxKf+/qlhMq02MUXppub3Kh4AAQCiAAAE6AW6AAsAlUAVBgUeCAgHBwADBB4CAQIKCR4LAAgHuP/AQB0QEjQHVANKIAogDQIKGg0ECSABIAABACAQEAJVALj/9rQPDwJVALj/9rQNDQJVALj/+rQMDAJVALj/+rQMDAZVALj/8EAKDQ0GVQBdDDtbGCtOEPQrKysrKytdPE39PE4Q9l1N9OQrAD88/Tw/PP08EjkvPBD9PDEwMxEhFSERIRUhESEVogQk/J4DK/zVA4QFuq3+P6z+Da0AAAEAqAAABIUFugAJAI1AKwYFHggIjwcBBwcAAwQeAgECAAgHnCACIAsCAhoLBAkgASAAAQAgEBACVQC4//a0Dw8CVQC4//a0DQ0CVQC4//pACwwMAlUADAsLBlUAuP/+tAwMBlUAuP/wQAoNDQZVAF0KO1wYK04Q9CsrKysrKytdPE39PE4Q9l1N5AA/Pzz9PBI5L108EP08MTAzESEVIREhFSERqAPd/OUCsP1QBbqt/jqt/WYAAQBt/+cFuQXTACUBE0AaGxQbFQJgJwFeCBMBEgMkJAAhEhcCJQAeAgG4/8BAIAwMBlUBAQYXHg4DIR4GCQEBJiclJCADAyACICdgAgMCuP/ktA8PAlUCuP/ytA0NAlUCuP/atAwMAlUCuP/0QBsMDAZVAnKAJwEnHSYgCgEKEAwMBlUKGSZjWxgrThD0K11N7U0QXfYrKysrXTxNEP08ERI5LwA/7T/tEjkvKzz9PBESORESOQEREjkSOTEwQ3lARAQjGxwaHBkcAwYMJhAlFSYfJgglBCYjJRgNHSEAFg8TIQEREhQTIAcdIQAiBSUhARwLFyEBFBEXIQEeCSEhACQDISEAACsrKysBKysQPBA8KysrKysrKysrKoEBXQBdATUlEQYEIyIkAjU0EiQzMgQWFwcuAiMiBgYHBhUUEgQzMjY3EQNMAm2P/tCg2P6ftLMBUNufAQGSJq8hYrZvhcJ3ITiHAQKRfvA+Aj+sAf3gcnO5AV7Y1gFztGe4lDBwgE1RhE+In8T++IBhNwERAAEApAAABSIFugALANi5AA3/wEAaExU0BAMeCQqgCtAKAgoFAgILCAgFCCAHBwa4/+60Dw8CVQa4//JACw0NAlUGEAwMAlUGuP/gQBgLCwZVBgEMDAZVBl2ADQENAgsgASAAAQC4/8BAChMVNAAgEBACVQC4//a0Dw8CVQC4//a0DQ0CVQC4//pACwwMAlUACAsLBlUAuP/3tAwMBlUAuP/4QBYNDQZVAF0MIA0BIA1QDWANcA0EO1kYK11xEPYrKysrKysrK108/TwQXfYrKysrKzwQ/TwAPzw/PDldLzz9PDEwASszETMRIREzESMRIRGkwgL6wsL9BgW6/aYCWvpGArP9TQABAL8AAAGBBboAAwDMtQECAAgCBbj/wLM4PTQFuP/AszM0NAW4/8CzLTA0Bbj/wLMoKTQFuP/AsyMlNAW4/8CzHR40Bbj/wLMYGjQFuP/AQCoNEDQgBZAFrwUDAyABAACPAKAAsAAELwBAAFAA3wDwAAUSIACPAJAAAwW4/8BACw0NAlUAGBAQAlUAuP/stA8PAlUAuP/utA0NAlUAuP/2QBAMDAJVACALCwZVAKIE1lkYKxD2KysrKysrXUNcWLKAAAEBXVlxcjz9XSsrKysrKysrPAA/PzEwMxEzEb/CBbr6RgABADf/5wNhBboAEQCpQBBlAmcGdAJ1BogNiBEGCQIBuP/AtAsMBlUBuAEaQAsEHg8JCSYKCggmC7j/6rQQEAJVC7j/6rQNDQJVC7j//rQMDAJVC7j/6LQLCwZVC7j//kAWDAwGVQtdIBMBIBNAE1ATYBMEEwEmALj/6LQMDAJVALj/6rQMDAZVALj/3EAKDQ0GVQBLErZZGCsQ9isrK+0QXXH2KysrKyvtPBDtAD/t7Ss/MTAAXRM3FhYzMjY2NREzERQGBiMiJjuvB3BjSWoowlnBgsHNAaAYqHxDc34D8vwZuMpq3gAAAQCWAAAFUgW6AAsB/kAeAyI3OQgJOicKNQY2CkcKVwOGA9cDB3YK2QPZCgMGuP/0QBgNDQJVKAWMBIoFqgTqCAUKBAE1BNYEAgm4/+BACRIhNAMgEiE0A7j/3rMMORIJuP/gsxIhNAi4/+CzEiE0BLj/4LMdITQEuP/AsxIWNAi4/95APRk5CAklJT0ICRkZPQYGBwkKCQgKBQMEBCAFChQFBQoJCAggBwYUBwcGCgoABQIEAQIHCwgACAoDAgsBAAS4AjpADzAFAaAFsAXABeAFBAVKCLgCOkALMAcBIAeAB7AHAwe4AoZADAsgIAABACAQEAJVALj/9rQPDwJVALj/9rQNDQJVALj/+rQMDAJVALj/+rQMDAZVALj/8kAKDQ0GVQBdDDuoGCsQ9CsrKysrK13t/V1x7fRdce0QPBA8PDwAPzw8PD88PDwSOS+HBS4rDn0QxIcFLhgrBH0QxAcIEDwIPAFLsBhTS7AbUVpYuQAE/9g4WbEGAkNUWLkABP/wswwRNAO4//BAFwwRNAYQDhE0CBAOEDQJEA4RNAoQDRA0ACsrKysrK1kxMAErKysrKysrQ1xYQBEJIhk5CCwZOQQsGTkEIhs5Bbj/3rYWOQQiFjkGuP/eQAsSOQgiFDkEQBQ5CLj/3rUlOQRAFTkrKysrKysrKysrK1kAKysrAXFyXSsAcV0rKzMRMxEBIQEBIQEHEZbCAtgBB/2ZAoL/AP328AW6/SkC1/2u/JgC5ur+BAABAJYAAAQqBboABQBtQAwBAgQDHgUACCAEAQS4AqdADwcCAyABIAABACAQEAJVALj/9rQPDwJVALj/9rQNDQJVALj/+rQMDAJVALj/9rQMDAZVALj/+EAKDQ0GVQBdBjtcGCsQ9isrKysrK108/TwQ5l0APzz9PD8xMDMRMxEhFZbCAtIFuvrzrQABAJgAAAYPBboAEALksQICQ1RYuQAI//ZACwwMAlUIDg0RAlUCuP/utA0RAlUFuP/uQCgNEQJVDBIMDAJVBQ8MAwkAAQIICQsOAAgJAgoLBhAQAlULEA0NAlULuP/6tgwMAlULEAC4/+a0EBACVQC4//i0Dw8CVQC4//y0DQ0CVQAvKysrzS8rKyvNAD8/wMAQ0NDAERIXOSsrMTABKysrABuxBgJDVFhAHwcgCwsGVQYgCwsGVQMgCwsGVQQgCwsGVQUgCwsGVQi4//JAIwsLBlUCDAsLBlUDBgwMBlUCDgwMBlUJDAwMBlUKDAwMBlUHuP/4tA0NBlUIuP/4QB8NDQZVJgUBDCAKEjQPIAoSNA8FDAMAAQ4LAAgIAQIKuP/utAsLBlUKuP/utAwMBlUKuwJWABIAEAJWQA0ADAsLBlUABgwMBlUAuP/4tA0NBlUAAS8rKyv0L/QrKwA/PD88PBESFzkrK10xMAErKysrKysrKwArKysrKxtAfwACDwgUAhsIBHYMhgzIDAMJDEkMSQ8DKQQlDSwOWANbBHYNeA6HDQgLAgUIOQ02Dk8CSwNEB0AITQ1CDgqYApkDlgeWCKgDpwcGEgIPDg4wBQIUBQUCCAwNDTAFCBQFBQgMUg9SAUABAgIICAkKCwsNDQ4OEAAICQJgEoASAhK6AqgADQExsgUgCLgBMUAKDAkKIEAMfwsBC7oCVgAOAQuyBSACuAELQAkPAQAgD3AQARC4Ala3IAVgBYAFAwW4AqizETtZGCsZEPRd9F08GP08EO0aGRDt9F08Ghj9PBDtGhkQ7eRdABg/Pzw8EDwQPBA8EDwQPBA8GhDt7YcFLiuHfcSHLhgrh33EMTAAS7ALU0uwHlFaWL0ADP/7AAj/1gAC/9Y4ODhZAUuwDFNLsChRWli5AA3/+LEOCjg4WQFDXFi5AA3/1LYhOQ4sITkNuP/Utjc5DjI3OQ24/9S1LTkOLC05KysrKysrWXJxXQBxXQFdWVkzESEBFhc2NwEhESMRASMBEZgBJAFbMBYZNQFfAQW7/lav/lgFuvvykUhQmwP8+kYEy/s1BOD7IAABAJwAAAUfBboACQF9sRILuP/AQAoTFTQIGAwWAlUDuP/oQCEMFgJVCAIDAyAHCBQHBwgCBwMDCAkEAgIJBwgEAyAGBgW4/+y0Dw8CVQW4//JACw0NAlUFEgwMAlUFuP/3QBoLCwZVBV0gCwEgC1ALYAtwC4ALBQsICSABALj/wEANExU0IAABACAQEAJVALj/9rQPDwJVALj/9rQNDQJVALj/+kALDAwCVQAECwsGVQC4//e0DAwGVQC4//hACg0NBlUAXQo7WRgrEPYrKysrKysrXSs8/TwQXXH0KysrKzwQ/TwAPzw/PBI5OQEROTmHBC4rh33EsQYCQ1RYuQAD/+C3DBE0CCAMETQAKytZMTArKwErQ1xYtAhARjkDuP/AtkY5CEAyOQO4/8C2MjkHIhk5Arj/3rYZOQciMjkCuP/etjI5ByIjOQK4/95ACyM5Bw4UOQcOEzkCuP/0thM5Bw4dOQK4//S2HTkHDhU5Arj/+LEVOSsrKysrKysBKysrKysrACsrKytZMxEzAREzESMBEZzHAwK6x/z+Bbr7gQR/+kYEgPuAAAACAGP/5wXdBdQADgAbAMpAUBoPARQQFBQbFxsbBAQQBBQLFwsbBKkXtg7GDgMXFxgbAiAdQBFPE08XQBpYBVgJVxBVEV8TWhdfGFYaVxuLF5kCEBkeAwMSHgsJFSYgBwEHuP/otBAQAlUHuP/utA0NAlUHuP/wtAwMAlUHuP/qtAsLBlUHuP/0tA0NBlUHuP/6QCEMDAZVBxqAHQEdDyYgAAEABgsLBlUABgwMBlUAGRxjXBgrThD0KytdTe1OEF32KysrKysrXU3tAD/tP+0xMAFdcQBdXV1xExAAITIEEhUUAgQjIiQCNxAAMzIAETQCJiMiAGMBiAE2ywFGq7T+tr/P/rqoyAEd19sBG3npkc7+1wLKAW0BncL+pdzf/qC1yAFavv73/s8BNAEbswELk/7lAAIAngAABP0FugANABgAskAsZRFrFAJLEEsUWxBbFAQLDB4PDg4AFxgeAgECAAgSJggKDQ0CVQgQCwsGVQi4//RAGwwMBlUIGiAaASAaARoYDSABIAABACAQEAJVALj/9rQPDwJVALj/9rQNDQJVALj/+kALDAwCVQAMCwsGVQC4//q0DAwGVQC4//BACg0NBlUAXRk7XBgrEPYrKysrKysrXTz9PE4QcV32KysrTe0APz88/TwSOS88/TwxMAFdAF0zESEyFx4CFRQCISERESEyNjU0JicmIyGeAimSTWySWe7+yf6IAXu8nl1MMYT+iQW6DhJltm27/v39rAMBjH9cgxUNAAACAFj/jgXuBdQAFQAoAWhAlV8mnyYCGRg3FQILHAQfBCMbHBQfFCMGKgUtFysmOwU8FzomTAVMF0kmXQVVI1gmbwV7A3oFjAOMBZUAmgOkAKsD1QDVFuUA5RflGBocBSsAKgU7BQRdBZIYlibVJgQlFiomNBY5JkkYSRxFH0UjSyZWCFgRVRVaHFodVh9XIFciaQVmFWsmeyaOHI4m2xjcJhkLGAEVuP/Ushs5ALj/1EA4GzkEGBQYKgU6BQQCAxYoAwcoJhgWBQAGIQMTGgUCKCYYFgAFJB4eDwMCCCQeBwkaJhMYDw8CVRO4/+60DQ0CVRO4/+i0DAwCVRO4//C0CwsGVRO4//S0DQ0GVRO4//RAJQwMBlUTSgIaICqAKgIqISYgCwELGAsLBlULBgwMBlULGSljXBgrThD0KytdTe1OEF32TfQrKysrKyvtAD/tPz/tERc5EjkBERI5Ehc5ABEzEMkQyV0xMAErK11dAHJxXQFdcXIlFhcHJicGIyIkAjU0EiQzMgQSFRQCJRYXNhE0AiYjIgAREAAzMjcmJwT1h3I5np2jxcf+vK+wAUXJywFGq2795qhtq3npkdn+4gEb3GhcW2WdXSuHOXtbwAFc2tkBZLrB/qXatf7fjS9dnAE5sgEKk/7X/tn+4v7OJzsZAAIAoQAABa0FugAYACIB/EAhEgsOARI2HFofZghtHwQJEA0NBlUIEA0NBlUHEA0NBlUkuP/AtAwMAlUNuP/0tAwMAlUMuP/0tAwMAlULuP/0tAwMAlUSuP/isxIaNBK4//CzIic0Ebj/4rMdJzQQuP/isx0nNA+4/+KzHSc0Erj/2LMdJjQRuP/isxIaNBC4/+KzEho0D7j/4kBJEho0JQ5KHEogUwtcHG0ccgl4DnkPhQqID5cNqQ+4D+gO5w8QDgwMIBEPFBERDxEPDAkSGwIhGhYKBhIREA0MBRgJCRYXGhkeF7j/wEAZCwsGVRcXACEiHgIBAgAYGA8PDggeJg6cBrj/6LQPDwJVBrj/9rQNDQJVBrj/4EAiDAwCVQYGDQ0GVQZdICRwJIAkAyQiGCABIAABACAQEAJVALj/9rQPDwJVALj/9rQNDQJVALj/+kALDAwCVQAGCwsGVQC4//e0DAwGVQC4//hACg0NBlUAXSM7qBgrThD0KysrKysrK108Tf08EF32KysrKxnkGO0APzwQPBA8Pzz9PBI5Lyv9PBA8OS8SFzkBERc5hw4uKwV9EMQxMAFdKysrKysrKysrKysrKwArKytdQ1xYQAoIQA85DxA6ERI6KysrWQFxQ1xYuQAO/95AGhk5ESIZORIiGTkOQBw5ECIUORAiHzkQIhU5KysrKysrK1kzESEyFhYVFAYHFhcWFxMjAy4CJyYjIxERITI2NjU0JiMhoQKKxMx6ytNNKFVM//TCVW5XLSFL4QGhhZZOl6P+MAW6T8h5nNYdJSROdf5xATGEjDgLB/11AzM3eUdohgAAAQBc/+cE6wXTADACFUAnYwNjBHMDdAQEJSc1AzkcQwNJB0wdRR9EJEYnUwNZB1wdVyiJEw4juP/ytBAQAlUkuP/ytBAQAlUluP/ytBAQAlUmuP/ytBAQAlUnuP/ytBAQAlUjuP/2tA0QAlUkuP/2tA0QAlUluP/2tA0QAlUmuP/2tA0QAlUnuP/2QEYNEAJVKA0mJAIkAyclNg80I0QlRS9aIFYjVSVsC2oNaw5mFGUYeQt6DXoPfRB1JHMlhgOKC4kNig+NEIUkgyWSDZYPlhUesQYCQ1RYQC0hJhIbJhoJJikBJgAAKRoSBDIxJgBlAAIADS15G4kbAhslFg0tHiclASUFFgW4//RADAwMBlUFHi0JHh4WAwA/7T/tKxESOV0REjkREjldERI5XQEREhc5L+0v7S/tL+0bQC0lJA4NCwUhHB0eGwgHBgQDAgYBJSQiDg0LBgUeGy0aQAwMAlWPGgEa7RYALQG4/8BAEgwMAlUQASABUAFgAXABkAEGAbgBsEATLR4eFgMFHi0JGyYaSgkmACkBKbj/6rQODgJVKbj/9EANDAwCVSkaMiEmEgEmErj/7LQODgJVErj/9rQNDQJVErj/+EAPDAwCVRJUIAABABkxY1sYK04Q9F1N5CsrK+0Q7U4Q9isrXU3t9O0AP+0/7RD9XSvkEP1dK/QREhc5ERc5ERI5OQESFzlZMTAAXXErKysrKysrKysrAV1xEzceAjMyNjY1NCYnJiQnJiY1NDY2MzIWFhcHJiYjIgYVFBcWBBcWFhUUBgYjIiQmXLcNX8h9b6pTUFw7/mxRaWd+8pSj+YYFug+tqbChOTgB2ViAeob7ncf+85kB1xBujVdCc0RFZyMXYSs3o2VvwWRpzIEOi46BW08zM2soO7V2dc9zdOkAAAEAMAAABLoFugAHAIlADQUCHgQDAgAIBwYFBAm4AnOzIAQBBLgBAbcGIAECLwMBA7gBAbUBASAAAQC4/+hACxAQAlUACA8PAlUAuP/ytAwMAlUAuP/itA0NAlUAuP/8tAwMBlUAuP/+tA0NBlUAuAJzswi2mRgrEPYrKysrKytdPBD0XTwQ/eRd5hA8EDwAPz88/TwxMCERITUhFSERAhP+HQSK/hsFDa2t+vMAAAEAof/nBSIFugAUANlACiYPWARYCMkIBBa4/8BAFhMVNDQEOwhGBEoIdg+mBegPBwwAAhG4Aru0BgkUJgK4/+y0Dw8CVQK4//JACw0NAlUCEAwMAlUCuP/gQBwLCwZVAl0gFgEgFlAWAmAWcBaAFgMWDSYgCgEKuP/AQAoTFTQKIBAQAlUKuP/2tA8PAlUKuP/2tA0NAlUKuP/6QAsMDAJVCgQLCwZVCrj/97QMDAZVCrj/+EAKDQ0GVQpdFTtZGCtOEPQrKysrKysrK13tTRBdXXH2KysrK03tAD/tPzwxMAFdKwBdATMRFAIEIyIkAjURMxEUFhYzMjYRBGDCZP771M7++nDCR6191rYFuvyx3f78o44BDekDT/yyv7ViwgEUAAABAAkAAAVGBboACgE+sQICQ1RYQBIFAQAIAgECAAgKAAUJCAUBAgUv3c0Q3c0RMzMAPz8/ERI5MTAbQCQvBQEqACgDJQovDDAMYAyJCIkJkAzADPAMCyAMUAwCBAILCAKxBgJDVFi3CQEMCwAIAQIAPz8BERI5ORtAJAoJCSAIBRQICAUAAQEgAgUUAgIFCQECBekgCgAICWUIAWUCCLj/wEALKDlQCAGACJAIAgi4AQFADQJAKDlfAgGPAp8CAgK4AQFAESAFUAUCMAVgBZAFwAXwBQUFuAKIswtgqBgrGRD0XXHkXXEr5F1xKxgQ7RDtAD88GhntGD88hwUuK30QxIcuGCt9EMQBS7ALU0uwFFFaWLIADwq4//GyCRIBuP/xsggUArj/7jg4ODg4OFkBS7AoU0uwNlFaWLkAAP/AOFlZMTABXXFdAF1ZIQEzARYXNjcBMwECQf3I0gF9Lh8iLQGMxv3CBbr714BweHgEKfpGAAABABkAAAd2BboAGAHbQCYpACYRKRImGDkANhE5EjYYSQBHEUkSRxhYAFcRWBJXGBCYCJgPArEGAkNUWEAzEAEaGSsVNAU0DEQFRAxLFVQFVAxbFWQFZAxrFXQFdAx7FQ8FFQwDAAESCAAIDwIIAgECAD8/Pz8/ERIXOV0BERI5ORtAHgMEBQUCBgcICAUKCwwMCQ0ODw8MFBMSEhUWFxgYFbj/PLMFABgguP88swwSESC4/zxAWhUICSAABQICIAEAFAEBABgFCAgeFRgUFRUYEgwJCR4VEhQVFRIRDA8PIBARFBAQERIJDAgYFQUPERAMAAIFFQwFAxgQDw8JCQgIAgIBAhgSEhERAAgaFxcaEEEJAVEAIAAMAVEAFQFRAEAABQFRtiAgAQEBGRm4AYuxqBgrThD0XRoZTf0aGP39Ghn9GE5FZUTmAD88EDwQPD88EDwQPBA8EDwSFzkBEjk5ERI5ORESOTkROTmHTS4rh33Ehy4YK4d9xIcuGCuHfcSHLhgrh33EKysrhw4QxMSHDhA8xIcOEMTEhw4QxMSHDhDExIcOEMTEAUuwD1NLsBFRWliyEgoYuP/2ODhZAUuwJVNLsCpRWli5AAD/wDhZAEuwC1NLsA5RWlizDEAFQDg4WVkxMAFyXSEBMxMWFzY3ATMTEhc2NxMzASMBJicGBwEBnv57x98kGjgKARfq0k8jHC3mw/5uu/7LJwcXFP7JBbr8P5eV6yQD3v0a/uzzi7QDrvpGBF2MIGVH+6MAAQAJAAAFSQW6ABMCtUApJhIBGQEWCwIpEikTOAE3AzgIOAk4DToONRI3EwoSEyASITQSIBIhNA64/+CzEiE0Dbj/4LMSITQJuP/gsxIhNAi4/+BAbBIhNAQgEiE0AyASITR3AXcLAiYEKQcoCyoOJhI2BDoIOgs6DjUSSAhUBF0IXAtaDlQSZwFlBGoIawtpDmUSdQR6CHkLeg13EncThgSKB4oKlQS4CLcSxgTJCNcE2AjZDtYS5wToCOgO5hIsBrj/6kARDBECVRAWDBECVQsIDBECVQG4//izDBECVbEGAkNUWEALDAAVFBAYChEGVQa4/+hADgoRBlUQBgACDQAICgICAD88PzwREjk5KysBERI5ORtAXQYHCAkJAQYFBAMDCxAQEw8ODQ0BEBANERITEwsBAAkCDQsDDBMKCwEGEAITCQoTEyAACRQAAAkDAg0NIAwDFAwMAwoJCQMDAgITDQ0MDAAILxUBFRcXGiAMQAwCDLgBX7cgCpAKwAoDCrgBuLVfAp8CAgK4AbhACga0QBBQEM8QAxC4AV9ACiAAGRQVwiFgqBgrK070GhlN/V0Y5RntXe1d/V0YTkVlROZdAD88EDwQPD88EDwQPIcFTS4rh33Ehy4YK4d9xAAREjk5OTkPD4cOEDw8CMSHDhA8PAjEhw4QPDzEhw4QxMTEWSsrACsrMTABXQBdASsrKysrKysrQ1xYuQAL/95ACxk5ASIZOQ4YGzkSuP/eshs5E7j/3rIbOQS4/+i2GzkIIhs5Cbj/wLIcOQ24/8BAHxw5E0AcOQNAHDkNDhYXPBMSFhc9CAkWFzwDBBYXPQu4/95ALhI5ASISOQsMHSE9AQAdITwLCh0hPQECHSE8CwwTFz0BABMXPAsKExc9AQITFzwrKysrKysrKysrKysrKwErKysrKysrKysrK1kBcQFdcTMBATMBFhc2NwEzAQEjASYnBgcBCQI3/gznAQpTIzFDASfT/f0CK/D+jx8hMRX+kAL8Ar7+iHU/UFcBhf1N/PkCCy01UB7+AQAAAQAGAAAFRgW6AAwBarYICToDBDsJuP/nsxIXNAi4/+dADhIXNAQZEhc0AxkSFzQJuP/YsxghNAi4/9hAOxghNAQoGCE0EiYEKQgqCi8OBGgBaAZoC94GBAUEAwMGCAcJBgYJBgMJCgwQAlUJIAoLFAoKCwYDBgkDuP/2QBYMEAJVAyACARQCAgEGDAsGAQMCAAELuAIZQAkKCgkDAgIACA64AhhACQwJUkAKgAoCCrgBtUANCwsMIAADUk8CjwICArgBtUAJAQEAFBAQAlUAuP/2QAsPDwJVAAwNDQJVALj/4rQMDAJVALgCGLYNDsIhYKgYKyv2KysrKzwQ9F3tEP08EPRd7RDmAD8/PDw8EPQ8ERIXOQESOYcuKysIfRDEBYcuGCsrCH0QxIcOxMSHEA7ExEuwF1NLsBxRWli0CAwJDAS6//QAA//0ATg4ODhZMTAAXQFdQ1xYQAkJIhk5CCIZOQS4/96xGTkrKytZKysrKysrKysrIREBMwEWFzY3ATMBEQI7/cvsASFQRUJeARzi/bcCbQNN/kZ8fHOQAa/8s/2TAAAB/+H+aQSK/usAAwAaQAwBPwACGgUAGQRDQRgrThDkEOYAL03tMTADNSEVHwSp/mmCggAAAgBK/+gEHAQ+ACgANwItQCwJDQkqGQ0aKikNKio5DTYVNxs6KkkqXQ1dKmoNaSpgMIoNhimaFpsaqQ0VKLj/6LQLCwZVJ7j/6EAZCwsGVaYZqii2GbsoxBnPKNIV3SgIRBYBHrj/9EARDAwGVRISDAwGVQUMDAwGVTW4/+BAVQwMBlUfFx8YKywqNDkEOSxJBEgsVghZK2YIaSt2DIcMyQz5DfkrETc0DgEEEC8kNBcyIRQYXylvKQIpHC8OPw6PDp8O/w4Fnw6vDu8OAw4MDw8CVQ64/+q0EBACVQ64//RAFRAQBlUODA0NBlUOBg8PBlUODhwDF7gCqrYYlRQcHAcAuP/0QBoMDAZVAEUnCjIcAwspYRBhAAYNDQJVACUhJLj/7LQQEAJVJLj/7EALDQ0CVSQEDAwCVSS4/+S0CwsCVSS4//S0CwsGVSS4/9xACxAQBlUkBg8PBlUkuP/8tAwMBlUkuAJbQA4nQAAmECYgJjAmryYFObj/wLQODgJVJrj/1rYODgJVJjE5uP/AQA0eIzQwOcA5AqA5ATkXuP/0QEEQEAZVFyUYIi8kvwbPBgIfBj8GAgYODw8CVQYMDQ0CVQYYDAwCVQYMCwsCVQYMCwsGVQYODQ0GVQYQDAwGVQYxOBD2KysrKysrK11x7fTtKxBdcSv2Kytd7fQrKysrKysrKzz9K+XlAD/tP+QrP+395BESOS8rKysrK11x7XEREjkREjk5ARESFzkxMABdKysrKwFxXSsrAHElBgYjIiY1NDY2NzY3Njc2NTQnJiMiBgcnPgIzMhYWFxYVFRQWFyMmAwYHDgIVFBYzMjY3NjUDPGS5aq+8R3NINWvaZwEzRYh/eR2wGG7QiYiqUBAJFyK8HBdixG9cMm1paKImHYNVRquFToFOFA4NGiQlCm4tPVlxGHGLS0BhSi548PuFPTgB3SgcEChNL0hgW089dwACAIb/6AQfBboAEAAdAYBAmwEFDA8kBTUFRQUFPx+wHwIfHyIcMxxCHHAfkB8GOhM8FjwaTBZMGl0IXQ1YD10WXhpqCGwNaA9uFm4awB/ZDNoX2hniE+wX7BnjHeAf/x8ZIAUvDy8UMAU/D0AFTA9QBWYF2h31BPoQDBAVDgQGAgAbHAYHAQoVHA4LGCTQCwEQC0ALYAuACwQfQA0NAlULDA8PAlULGA0NAlULuP/2tAwMAlULuP/wtAsLBlULuP/0tA8PBlULuP/gtAwMBlULuP/0QC8NDQZVC3QBETMABAwMAlUABA0NBlUAMwMlAgLAAQGQAaABsAHwAQQfAT8BTwEDAbj//rQQEAJVAbj//EAdDg4CVQEMDQ0CVQEQDAwCVQESCwsCVQEMCwsGVQG4//i0EBAGVQG4//xAFg8PBlUBGAwMBlUBFA0NBlUBGR5HNxgrThD0KysrKysrKysrK11xcjxNEP30KyvkEP0rKysrKysrK11x7QA/7T8/7T8RORESOTEwAF0BXXFyAHEhIxEzETYzMh4CFRAAIyInAxQXFjMyNjU0JiMiBgEtp7RysWKvcUD+8r28awI0VZF2rKV1dqwFuv31j0+PynP+7/7WnQGWv1WLzcvQxs0AAQBQ/+gD7QQ+ABoBWrECAkNUWEA0Dn8PAQ8LAUAAUABwAAMABBIcCwcYHAQLAQ4VBwgODgJVBwwNDQJVBwwMDAJVBxALCwJVBy8rKysrzdTGAD/tP+0QxF0yEMRdMjEwG0BHCQwBHxxDE0MXUxNTF2ATYBebApsDmg2kEKQaDAgNGQpqAmkDagV1DHANgA2mDLUJtgq1DAwWDIYM4wIDDiJfD28Pfw8DDwG4AqpAeTAAQABQAGAAcACQAKAA4ADwAAkADw8LAAAEEhwLBxgcBAscDwEPJA4IDQ0GVQ4iGwABACQLKx8BAQABAQFACwsGVQFAEBAGVQFIDAwGVQEaDQ0GVQFJHBUkzwcBHwc/BwIHDgsLBlUHChAQBlUHEgwMBlUHMRs0xBgrEPYrKytdce0Q9isrKytdcktTI0tRWli5AAH/wDhZ7XL0K+1yAD/tP+0SOS8ROS8QXeQQXeQxMABdcQFdcVkBFwYGIyIAETQSNjMyFhcHJiYjIgYVFBYzMjYDPLEd767a/vdy6Ymt3B+vGX9aiKqkhGqOAYUXt88BHQEKrAECga+hG2tsw9PWwoIAAAIARv/oA98FugARAB0BVUCkCgIEDSUNNA1EDQU1FDUcVwJUClIUUxxnAmQFZQljFGAcwB/UBdUT3RnlE+UU7xfrGeUd4B//HxYfHysaPBY8GksacB+QHwcuAiQNLhY6AjUNSwJFDUYUSRxXClYNZw3lBucW+gH0DhABFQMOCxAPABscCwcRAAoVHAMLGDMBACURDyUQENARARARQBFgEYARBB9ACwsCVR9ADQ0CVRESEBACVRG4//RAEQ8PAlURBg4OAlURGA0NAlURuP/yQAsLCwZVEQ4QEAZVEbj/7rQMDAZVEbj/+EBCDQ0GVRF0EiS/B88H3wf/BwQfBz8HTwcDBx4LCwJVBxgMDAJVBx4NDQJVBwwLCwZVBwwNDQZVBxoMDAZVBxkeNFAYK04Q9CsrKysrK11xTe39KysrKysrKysrK11xPBDtEP085AA/7T88P+0/PBE5ERI5MTAAXQFxXQBxITUGIyImJjU0EjYzMhYXETMRARQWMzI2NTQmIyIGAzhlxH/VdWrUg2CWL7P9IKx1dqWoe3ihhp6M+6OfAQOKUUECDvpGAhLMysHG2szEAAACAEv/6AQeBD4AFQAdAVNAFx8AHBUCVQNdBV0JVQtlA2sFbwllCwgVuP/ktA0NBlURuP/kQFINDQZVHRwNDQZVJxLZBfoU9hoEMRI6GTEcQRJNGkEcURJcGVIcYRJtGmEceAZ4FfYC9hgQABYBDw0XF1AWYBZwFgMWHA+QEKAQAhAQBBscCgcAugKqAAH/wLQQEAJVAbj/wEAQEBAGVRABAQGVExwECxdADbj/3LQNDQJVDbj/7rQNDQZVDbj/6rQMDAZVDbj/wEAJJyo0sA0BDRofuP/AsyUmNB+4/8BAQR4jNDAfAR8WMxAkB0AkKjQfBz8HTwcDByALCwJVBxgMDAJVBxwNDQJVBw4LCwZVBxwMDAZVBxYNDQZVBxkeNDcYK04Q9CsrKysrK10rTf3kThBxKyv2cSsrKytN7QA/7f1dKyvkP+0SOS9dPP1xPAEREjk5EjkxMAFdAF0rKysBcXIBFwYGIyIAERAAMzIAERQHIRYWMzI2ASEmJyYjIgYDXros7rnp/u8BFNzVAQ4B/OgKsoVjjP3aAlEMOFaJfKkBVhejtAEfAQMBDAEo/t7++RAgr7poAZWGQ2imAAEAEwAAAoAF0wAXAQ1AHhQJAQ8ZLxkwGUAZcBmbDJwNqQ0IGg0oDbAZwBkEGbj/wEAoGh80HQgNAwwPHAoBFQIrFBMEAwYACp8UART/E0AEFyUEAAMCkgEBALj/wLMxODQAuP/AQCscHzSQAAEZQA8PAlUZQA0OAlUAFBAQAlUAKA8PAlUAIg4OAlUALA0NAlUAuP/yQAsMDAJVABQLCwZVALj/6rQQEAZVALj/5rQPDwZVALj/+rcMDAZVAKMYGbwBugAhAPYBCgAYKyv2KysrKysrKysrKytdKys8EPQ8EDztEO3tXQA/Pzw8PP08P+05ETkxMEN5QBQQEQYJBwYIBgIGEAkSGwARBg8bASsBKyqBgQErcV0AcjMRIzUzNTQ3NjYzMhcHJiMiBhUVMxUjEbKfnxMag3ZMXBs4MlJEz88DmoxxazRGVxKdCkZgYoz8ZgACAEL+UQPqBD4AHgAqAW9AYAsLBRQsCyUUTAtFFAYJHRkdLAsmFCwjOQs2FEoLRhRWB1gLaAv6CvUVDi4jLCc+Iz4nTCeQLKAsBzYhNik/LEYLRiFFKVQhVClpB2MhYylgLIAs2ifoIe4j7ycRFxYGFbgCsbQoHBMHAbgCqkAQIAAwAGAAcACAAMAA0AAHALgCfUAyBRwcDwpFIhwMChYVMyUzCiUYGNAXARAXQBdgF4AXBCxACwwCVSxADQ0CVRcSEBACVRe4//RAEQ8PAlUXBg4OAlUXFg0NAlUXuP/qQAsLCwZVFxIQEAZVF7j/7rQMDAZVF7j//EBKDQ0GVRd0DwElACIfJL8Pzw/fD/8PBB8PPw9PDwMPIAsLAlUPGgwMAlUPIg0NAlUPHAsLBlUPDA0NBlUPGgwMBlUPGSssdCE0UBgrK070KysrKysrXXFN7fTtEP0rKysrKysrKysrXXE8EP3k9jwAP+3kP+39XeQ/7eQ/PDEwAV1xAF1xFxcWFxYzMjY3NicGIyICNTQSNjMyFzUzERQGBiMiJhMUFjMyNjU0JiMiBmavCzJDdH2IGA4BdrDb8G7Rjbx6pmXboL7qmaZ9fKitenioWBpRJTJkWjewiwE83ZgBAYyYgPxq+M94qwMq0cC/zMPGwwAAAQCHAAAD6AW6ABQBYbkAFv/AsxUXNAO4/+BADg0NBlUlBDUDRQO6DQQDuP/gQDoXGTQXCBEMERQDBQEADxwFBxQLCgwlCUAzNjT/CQHACQEWQAsLAlUWQBAQAlUJKBAQAlUJFA4OAlUJuP/sQBENDQJVCQQMDAJVCRoLCwJVCbj/9kALCwsGVQkUEBAGVQm4//hACw0NBlUJCg8PBlUJuP/2tgwMBlUJTha4/8BAFzQ2NLAW8BYCcBagFrAW/xYEFgIUJQEAuP/AQBAzNjTwAAEAACAA0ADgAAQAuP/6tBAQAlUAuP/6QBcODgJVAAQMDAJVAAgLCwJVAAQLCwZVALj/+kAWDw8GVQACDAwGVQACDQ0GVQBOFUdQGCsQ9isrKysrKysrXXErPP08EF1xK/QrKysrKysrKysrKytdcSvtAD88P+0/ETkROQESOTEwQ3lADgYOByUOBgwbAQ0IDxsBACsBKyuBACtdKwErMxEzETYzMhYWFREjETQmIyIGBhURh7R+wHauS7R1a1CNPAW6/fKSXaSc/V8CoYd7U459/bsAAgCIAAABPAW6AAMABwDNQF4JNgsLAlVPCZAJoAmwCcAJ3wnwCQcACR8JcAmACZ8JsAnACd8J4An/CQofCQEAAQcEAgMJBgN+AQAGBQYECgYHJQUABJ8EoASwBMAE4AQGwATwBAIABCAE0ATgBAQEuP/4tBAQAlUEuP/6QBcODgJVBAQMDAJVBAoLCwJVBBQLCwZVBLj/6rQQEAZVBLj//rQNDQZVBLj//EAKDAwGVQROCEdQGCsQ9isrKysrKysrXXFyPP08AD8/PD/tARESOTkREjk5MTABXXJxKxM1MxUDETMRiLS0tATrz8/7FQQm+9oAAAL/ov5RAToFugADABIA1UBFBAUlBTsEMwWGBQUXCAUFBwQEAgQFEwABDQsCAxQMBBEFCwcDfgEACwYHHBEPkBQBFBcXGgwMDSUKCpALAR8LPwtPCwMLuP/6QDcODgJVCxANDQJVCxAMDAJVCwwLCwJVCx4LCwZVCwwQEAZVCwgMDAZVCwwNDQZVCxkTFK0hR1AYKytO9CsrKysrKysrXXE8TRD9PE4QRWVE5nEAP03tPz/tERI5EjkBERI5ORESOTkRMzOHEAg8MTBDeUAOCBAPJggQChsBCQ4HGwAAKwErK4EBXRM1MxUBNxYzMjY1ETMRFAcGIyKGtP5oIjYfNza0M0GXSQTp0dH5e5kOSZIEXPugxE1kAAABAIgAAAP4BboACwJhQBsGDA0NBlUHBlYGWgkDDw3zBfYGAwkMEBACVQa4//S0DAwCVQq4//S0DAwCVQm4//S0DAwCVQO4/+hAEA0NBlVVA3cKAhIGIBMhNAi4//CzEic0Cbj/8LQSJzQSBbj/8LMSITQJuP/wQIQSJzQGBAQFBAY3CUcEBSUGLQpYCncDdQraA+MGB6YGASMGJgclCDkGOAk/DU8NWQRZBlgHWQl9BHkFmQnGBtIE1gbkBukH9wb5CBUSCgoFAwMEAgYGBwkJCAoKBQkICCUHBhQHBwYDBAQlBQoUBQUKCgkGAwQIAQIABAUGBwgICwsACgS4AQ9ACQUEDAwGVQUiCLgBD0AhIAc/BwIHEAwMBlUHGpANAQ0LJQACJQEBkAABPwBPAAIAuP/+QDEODgJVABANDQJVABAMDAJVAAoLCwJVABILCwZVABIMDAZVAAgNDQZVABkMDeEhR2YYKytO9CsrKysrKytdcTxNEO0Q7U4QcfYrXU3t9CvtAD88EDwQPD88PzwRFzmHBS4rBH0QxIcFLhgrDn0QxAcQCDwIPAMQCDwIPLEGAkNUWEANSwkBHwmEAwIJGA0RNAArXXFZMTABQ1xYQAoJLB05CQgdHTwGuP/esh05Brj/1LIgOQa4/9SxITkrKysrK1ldAHFdAXEAKytDXFi5AAb/wLIhOQO4/8CyFjkDuP/eshA5Brj/3rIQOQO4/96yDDkDuP/esQs5KysrKysrWQErKytDXFhAEt0EAQgUFjkJCBQUPAkIFBQ8Brj/9rIYOQa4/+yxGzkrKysrKwFdWQBdKysrKysBXXErMxEzEQEzAQEjAQcRiLQBqun+agG/3v6hfwW6/LwBsP52/WQCH3r+WwAAAQCDAAABNwW6AAMA47YFNgsLAlUFuP/Aszc4NAW4/8CzNDU0Bbj/wLMwMTQFuP/AsyIlNAW4/8BAJRUXNA8FHwWfBd8FBE8F3wXwBQMfBXAFgAX/BQQBAAAKAgMlAQC4/8CzNzg0ALj/wEAVMzU0nwABwADwAAIAACAA0ADgAAQAuP/4tBAQAlUAuP/6QB0ODgJVAAQMDAJVAAoLCwJVABQLCwZVAAgQEAZVALj//rQNDQZVALj//7QMDAZVALj//EAKDAwGVQBOBEdQGCsQ9isrKysrKysrK11xcisrPP08AD8/MTABXXFyKysrKysrMxEzEYO0Bbr6RgAAAQCHAAAGJgQ+ACMBx7kADf/0tA0NBlUIuP/0tA0NBlUJuP/YQE0LDTQlBOQE5AnhF+UgBdUF9iACFwggIwkYGyAJAwMjHhwGFRwLCwYHAQYjGhkQCtAlAZAloCUCJRcXGg4lkBEBEQQQEAJVERgPDwJVEbj/7EALDg4CVREUDAwCVRG4/+hAFwsLAlURAgsLBlURDBAQBlURBg8PBlURuP/6tAwMBlURuP/4tA0NBlURuAFdQAwYJZAbARsYDw8CVRu4/+xACw4OAlUbFAwMAlUbuP/uQBELCwJVGwQLCwZVGwoQEAZVG7j//kALDQ0GVRsMDw8GVRu4//y0DAwGVRu4AV1AFgACMyMlAdAAAZAAoAACHwA/AE8AAwC4//5AHQ4OAlUAEA0NAlUAEAwMAlUADAsLAlUAFgsLBlUAuP/8tBAQBlUAuP/0QBQPDwZVAAoMDAZVAA4NDQZVABkkJbgBeLMhR1AYKytO9CsrKysrKysrK11xcjxN/eQQ9CsrKysrKysrK13t9CsrKysrKysrKytd/U5FZUTmcXIAPzw8PD8/PE0Q7RDtERc5ARESORI5MTBDeUAODBQTJhQMERsBEg0VGwEAKwErK4EBXQBdKysrMxEzFTY2MzIWFzYzMhYVESMRNCYmIyIGFREjETQmIyIGBhURh6Eypmp2lx9+yp6qsyNcPnCUtFhkTIE6BCaVTl9iWLqvtv0nAp1sXzqVpP2XArJ4eFCakf3ZAAABAIcAAAPmBD4AFgF9QBMFAwYTAqgQuBDjA+cT8AP2EwYEuP/wQDwLDTR5EAGYENAY4Bj/GAQgCBQOFBYSHAUHAQYWDQoNDgwOJBhAEBACVRhACwsCVQsoEBACVQsUDg4CVQu4/+xAEQ0NAlULBAwMAlULIgsLAlULuP/0QAsLCwZVCxQQEAZVC7j/+UALDQ0GVQsKDw8GVQu4//ZAEgwMBlULQDM2NP8LAf8LAQtOGLj/wEAaNDY0sBjwGAJwGKAYsBjAGAQYAwIzFRYlAQC4//a0ERECVQC4//q0EBACVQC4//pAFw4OAlUABAwMAlUACgsLAlUABAsLBlUAuP/6QBEPDwZVAAIMDAZVAAQNDQZVALj/wEASMzY08AABAAAgANAA4AAEAE4XEPZdcSsrKysrKysrKys8/Tz0PBBdcSv2XXErKysrKysrKysrKysr7TwQPAA/PD8/7RE5ARI5MTBDeUAWBhEJCggKBwoDBhAmEQYOGwEPChIbAQArASsrKoEBXXEAK11xMxEzFTYzMhYWFxYVESMRNCYmIyIGFRGHonXdYKFQEAq0KmtIc6cEJpevRXBNMn39cwKGbm1Bksz9vAAAAgBE/+gEJwQ+AA0AGQFrthUYDQ0GVRO4/+i0DQ0GVQ+4/+hAcw0NBlUZGA0NBlUSBwoZDEcGSAhWBlkIZwZpCAg0EDoSOhY1GEUQSxJLFkUYXAVcCVIQXRJdFlIYbQVtCWQQbRJtFmQYdwEVCQYFDVsDVAVUClsMbANlBWUKbAwKFxwEBxEcCwsUJBtADQ0CVRtACwsCVQe4/+pAEQ8PAlUHGA0NAlUHEAsLAlUHuP/wtAsLBlUHuP/wtA0NBlUHuP/wtA8PBlUHuP/wtAwMBlUHuP/AQBMkJTQwBwEABxAHIAcDBzHfGwEbuP/AQEkeIzQwGwEbDiQADA4PAlUAEg0NAlUADAwMAlUAHAsLAlUADgsLBlUADg0NBlUADBAQBlUAFgwMBlUAQCQlNB8APwACADEaNDcYKxD2XSsrKysrKysrK+0QcStd9l1dKysrKysrKysrK+0AP+0/7TEwAXFdAHFDXFhACVMFUwliBWIJBAFdWQArKysrExA3NjMyABUUBgYjIgATFBYzMjY1NCYjIgZEpInF2wEWe+uL3/7tubKHhrKzhYeyAhMBJ452/uH9zeuCAR4BDczLzNHFy8oAAgCH/mkEIQQ+ABIAHgFiQI4MEC0QPRBLEAQ/ILAgAh8gKQwjHTIVMh1CHXAgkCAIOhc6G0oXShtZCFsMXBdcG2oIawxpEG0XaxvAINMU3RjdGtMe5BTkHuAg/yAWIwQrECsVNQQ6EEYEShBaEOUL6x3+EAsRDgMWHBwGBwEGFhwOCwAOGSTQCgEQCkAKYAqACgQgQAsLAlUgQA0NAlUKuP/mQAsPDwJVChgNDQJVCrj/+rQMDAJVCrj/7rQLCwZVCrj/9LQPDwZVCrj/6EAjDAwGVQp0ARMzAjMSJQAAwAEBkAGgAbAB8AEEHwE/AU8BAwG4//xAHQ4OAlUBEA0NAlUBEAwMAlUBEAsLAlUBDAsLBlUBuP/2tBAQBlUBuP/8QBYPDwZVAQwMDAZVARINDQZVARkfRzcYAStOEPQrKysrKysrKytdcXI8TRD99OQQ/SsrKysrKysrXXHtAD8/7T8/7RE5EjkxMABdAV1xcgBxExEzFTY2MzIWFhUUAgYjIiYnEQMUFjMyNjU0JiMiBoekOpJoiNBqdd97Wo8uEaZ2eKundHOx/mkFvYpRUYz/mKP++4tMOv37A6TNxMvVy8rXAAACAEj+aQPgBD4AEAAcATZAjgsCKwIqGDsCSwJ5DAY/FT8ZSxmQHqAeBTQTNBs/HkQTRBtTE1MbYxNjG2AegB7UBtUS5gbpDOoYECkCIgwrFTkCNQxJAkYMWgJpAtkM2xjjFukZ5hv8Ag8BBA0UGhwLBw4GFBwECwAOFw4zACUQENAPARAPQA9gD4APBB5ACwwCVR5ADQ0CVQ8SEBACVQ+4//RAEQ8PAlUPBg4OAlUPFg0NAlUPuP/+QAsMDAJVDxYQEAZVD7j/6LQMDAZVD7j/9EA/DQ0GVQ90ESS/B88H3wf/BwQfBz8HTwcDByQLCwJVBxoMDAJVByINDQJVBxYMDAZVBxoNDQZVBxkdHnQhNFAYKytO9CsrKysrXXFN7f0rKysrKysrKysrXXE8EP30PAA/P+0/P+0RORI5MTAAXQFdcQBxAREGBiMiABE0NjYzMhc1MxEBFBYzMjY1NCYjIgYDLCqXVb3+72/TfsVxov0hrHhzpq92daP+aQIIO04BLgEHoP6Dpo76QwOtzc3Dx9TWxwAAAQCFAAACxgQ+ABEAyUA7LxMBEAQBIwQ0BEMEUwRmBHQEBgkRCAkICQ0TEQkNAAMIAQscBgcBBgAKCSiQCAEIIiATARMCIhElAQC4/8BAEDM2NPAAAQAAIADQAOAABAC4//i0EBACVQC4//hAEQ4OAlUABAwMAlUABgsLAlUAuP/8tBAQBlUAuP/0QBYPDwZVAAYMDAZVAAgNDQZVAE4SR8QYKxD2KysrKysrKytdcSs8/eQQXfRy5AA/Pz/tETk5ETk5ARESOTkAEMmHDn3EMTAAXXIBXTMRMxU2NjMyFwcmIyIGBwYVEYWiPmk/W14+QkI7XhQeBCahcUg6pydHP2By/dQAAAEAP//oA7EEPgAwAxdAewQiFCI6CUoJRCRWImUifAmOCYQkphOrLMIDDQkXGhgXMEss1hcFGwJVAgIQMgEKGFwIXAlcClwLXAxcDWoIaglqCmoLagxqDbQmtCcPJyYkJyQpNiRaClkLZCZkKHQjdCSAJJMKnAySKJcslTCkCqkMoyekKLMmxSYWKLj/9LQNDQZVIrj/9LQNDQZVI7j/9LQNDQZVJLj/9LQNDQZVKLj/9LQMDAZVIrj/9LQMDAZVI7j/9LQMDAZVJLj/9LQMDAZVHbj/3kASHjlaCCclDAoEGiAmFQQLLh0auAKqQCIZLAsLAlUfGT8ZTxlfGa8ZzxkGDxkfGW8Z3xkEHxmPGQIZvQJVABUAAAKqAAH/wEAUCwsCVRABQAECEAHQAQIAARABAgG4/8CzFBY0Abj/wEAQDhE0AQEuXB1sHQIdHBUHBLj/9LQLCwJVBLj/5rQQEAZVBLj/5kATDw8GVQQcLgsfGgEaJBlAExg0Mrj/wEAvDw8CVRkYDw8CVRkYDQ0CVRkWDAwCVRkgEBAGVRkgDw8GVRkQDAwGVRkWDQ0GVRm4AluyByQquP/AtRw50CoBKrj/5rQMDAJVKrj/6LQPDwJVKrj/6LQMDAZVKrj/6rYNDQZVKhoyuP/AQCEnKjRgMsAyAj8ygDICMhABAQEkABgNDQJVABANDQZVACC4//S0DQ0CVSC4//S0EBAGVSC4//RAGQ8PBlUgJA8QCwsCVQ8WDAwCVQ8gDQ0CVQ+4//pAIA8PAlUPDgwMBlUPDA0NBlUPIt8AAT8ATwACABkxNDcYK04Q9F1xTfQrKysrKyvtKysrECsr7XJOEF1xK/YrKysrcStN7fQrKysrKysrKyvtcgA/7SsrKz/tcRI5LysrXXFyK+QQ/V1xcivkERI5ERI5ARESFzkxMEN5QEAnLR4jBRQsJhEQEhATEAMGIg0gGwAJKAcbAQUtBxsBHhQgGwAhDiMbACIjDQwIKQobASgnCQoGKwQbAB8QHRsBACsrEDwQPCsQPBA8KwErKysrKiuBgYEAKysrKysrKysrXXEBXXJxXRM3FhYzMjY1NCcmJy4CNTQ2NzY2MzIWFhcHJiYjIgYVFBcWFxYXHgIVFAYGIyImP7IPiXt8eDUlk8aZT0E4KpFTfb1aEbAMc2l8ahYWLxuEv5dWacZ9z9kBPRxrcmVEPSMYJTJJgU5HeSgfK0h7ZxhSXFI3IxwdEwokM0F8XFqfV6wAAAEAJP/yAioFmQAXANi5AAr/wLMjJjQJuP/AQEEjJjSAGQEAAQwNCgEDABYQCSsPCgYWHAMLDxAiACIBDRIlDAH/BwhFCUVgB3AHgAeQBwQAByAHoAewB8AH0AcGB7j/7rQQEAJVB7j/9LQPDwJVB7j/8rQODgJVB7j/+LQNDQJVB7j/+LQMDAJVB7j/+rQQEAZVB7j/8EALDw8GVQcGDAwGVQe4/+i0DQ0GVQe6AmoAGAE2sWYYKxD2KysrKysrKysrXXH05BDtPP08EOT0PAA/7T88/TwRORI5ETMzEMkxMAFdKyslFwYjIiYmNREjNTMRNxEzFSMRFBYWMzICEBpMPGJsLISEs7W1EysoHqGfED5logJjjAEHbP6NjP2TTSwaAAABAIP/6APgBCYAGAFPuQAa/8BACRUXNAIgExY0D7j/8EAzEhQ0KxMBJAgTFgwBExYLBgAKERwDCwAzFiUYF0AzNjQaQBAQAlUXKBAQAlUXEg4OAlUXuP/sQAsNDQJVFwQMDAJVF7j/9EALCwsGVRcUEBAGVRe4//hACw0NBlUXDA8PBlUXuP/2QA0MDAZV/xcBwBcBF04auP/AQBU0NjSwGvAaAnAaoBqwGv8aBBoMJQm4/8BAEDM2NPAJAQAJIAnQCeAJBAm4//i0EBACVQm4//hAEQ4OAlUJBAwMAlUJCgsLBlUJuP/2QBYPDwZVCQIMDAZVCQINDQZVCU4ZR1AYKxD2KysrKysrK11xK+0QXXEr9l1xKysrKysrKysrKys8/eQAP+0/Pzw5OQEREjkxMEN5QBoEEA4NDw0CBgcIBggFCAMGEAQMGwANCBEbAAArASsqKoEAXQErKyshNQYjIiYmJyY1ETMRFBcWFjMyNjY1ETMRAz981V6jTxALtAsRblFRjju0nLRIbU81cwKS/bONMUdRU4+IAjn72gABABoAAAPoBCYACgHqsQICQ1RYQBcFCAAKCAYBBgoABQkIBQECBSQPDwJVBS8r3c0Q3c0RMzMAPz8/EjkxMBu3NQUBACIROQq4/95ADRE5CRYSHDQIFhIcNAK4/+qzEhw0Abj/6rMSHDQKuP/YQAkeITQAKB4hNAq4/+hACSIlNAAWIiU0Crj/2kB+KC40ACAoLjQPDCkAKAkmCjkANQpIAEcKVgFWAlkIWAlmAWYCaQhpCXgAdwF3AnkIeAl3CocBhwKGA4kHiAiKCZ0AmAmRCqwAogq9ALcHsQrJAMUK2gDVCuwA4wr7APQKLAoABQoYABYKKAAmCjcKTwBACgkFQBIWNAVACw00sQYCQ1RYQAkFAQAIBgEGAAq4//RADw0NBlUKAAwNDQZVAAUJCLj/9EASDQ0GVQgFAQIMDQ0GVQIFBQwLERI5L90rzRDdK80QzSvNKwAvPz8REjkxMBtANwoHCAglCQoUCQkKAAMCAiUBABQBAQAFCgoACgkICAICAQYHCgkDAAEFLwwBDCIIQEBACYAJAgm4ARu1QAWABQIFuAEbQAkgAkABIgvq0hgrEPbtGhn9Xf1dGhjt5F0REjk5Ejk5AD88EDwQPD88ETmHBS4rh33Ehy4YK4d9xFkxMAArKwFxXSsrKysrKysrKysrKwBdWSEBMxMWFzY3EzMBAa7+bL7kJR8YK+y5/m4EJv2EZ29UdgKI+9oAAAEABgAABbcEJgASBB2xAgJDVFi5ABL/9EARDQ0CVQcGDQ0CVQAGDQ0CVQq4/9S0DA0CVQS4/+hACwwNAlURIAwNAlUKuP/AtA4QAlUEuP/AQC8OEAJVEUAOEAJVBAoRAwEADAYHBgEGDwoACg0MBgwMAlUMEQECBAoEEQoMDAJVEbj/+LQNDQJVES8rK83NENbNENQrzQA/Pz8/PxESFzkxMAArKysrKysBKysrG0AWDxQBKgQpCgJKEVsRjhEDESANDQZVCrj/4LQNDQZVBLj/4LQNDQZVEbj/8EAJHyE0EBwdJzQJuP/wQLcfJDQEBgwJEwYbCRkSBQQABAYLCQsOCBIQABMDFAccCBsLHQ4kACUHKggrDjQANQc6CDsORANHBkAHTQhLC0MPRxFKElsPUhJrB2QIZxJ5BnoHdAi5BroPthL1BvsJKAsRKAAoDScOKA8nEi8UOAA3EncIhgiYA5cMpwGoAqgLpgy1ALYGug7IBNYG2QnoBOgP5xL0BvoJHAsGDQ0GVQwGDQ0GVRAGDQ0GVQ4GDQ0GVQ8GDQ0GVRKxBgJDVFhAGwoODwQSABEIBwglBw8lDhIlAAAOBwMNAQwlDbj/1kA3CwsGVQ0CJQEqCwsGVQENARQTBgoLESYKKxFUBFIKXBFsEXwRihEKEQoEAwABDwoACgwGBwYBBgA/Pz8/PxESFzldARESOTkvK/QvK/QREhc5EOQQ5BDkERI5ERI5ERI5G0AUAwUFAgYHBwUJCgoICwwMChAREQ+4/0uzBQASILj/SUBmCg8OIMMRBwggBxESEisFBxQFBQcOCgwMJQ0OFA0NDggRDw8rCggUCgoIAAUCAiUBABQBAQAAAgEHEgQIDxEMDg0KEQoEAxINDAwICAcHAgIBBhIPDw4OAAoU9hANAWANcA2ADQMNuAGnQAogTwoBbwp/CgIKuAJVQAlPEQFvEX8RAhG4AlVACxAFAWAFcAWABQMFuAGntQH2E/ZmGCtOEPQZTfRdXRj9XXH9XXEaGf1dXRjmAD88EDwQPD88EDwQPBA8EDwSFzkBERI5ORI5ORE5ORI5OYdNLiuHfcSHLhgrh33Ehy4YK4d9xIcuGCuHfcQrKyuHDhDEBw4QPAcOEDyHDhDEhw4QxEuwH1NYtA0gDCACvP/gAAH/4AAO/9C0ADAPIBK4/+ABODg4ODg4ODhZS7A0U1i5AAj/0LEHMAE4OFlLsCFTS7AzUVpYuQAI/+CxByABODhZS7ASU0uwHlFaWLkADv/Qtg8gDSAMIAi4/9CyBzASuP/gsgA4Arr/4AAB/+ABODg4ODg4ODg4OFlLsBJTS7AXUVpYuQAR/+CzCiAEIAA4ODhZWTEwAUNcWLkADv/UthI5ACwSOQC4/9SxEzkrKytZKysrKytdcXIrKysAKysrcV0BXVkhATMTFzY3EzMTFzcTMwEjAycDAUv+u7qpPwQzqbmfNT22r/60u6kp1wQm/ZvkEcoCbv2Yy80CZvvaAny1/M8AAQAPAAAD8QQmABAB3LECAkNUWEAVDwELBgQCCQYCBg0KAAoPGA8PAlUPLysAPz8/PxEXOTEwG7cPEgEPIhk5Brj/3kBQGTlaD5YElgiZDpoPwAXABsAHyw8JD0AWORoDEwkVDRoQNQE6C4EBjgsILxJXBFkHWQtYDpcBmAqYC7cCuAzIC8oOzBDaA9UJ0Q3bEOUKEhKxBgJDVFhACwwAEhEPGA0QBlUGuP/oQA4NEAZVDwYAAg0ACgoCBgA/PD88ERI5OSsrARESOTkbQGYGBgMHCAkJAQYGCQUEAwMLDw8QDg0NAQ8PDRALAQAJAg0LAwwQCgYPAg8KEMYAxgkCECUACRQAAAkDAg3GDQENJQwDFAwMAwoJCQMDAgYQDQ0MDAAKTxIBEkkNfgwiCg9hBgl+QAq4ARu3QAZQBoAGAwa4AkNADiADfgIiTwABAEkRfMQYKxD2XfTtGhn9Xf0aGO0Q5RD07eZdAD88EDwQPD88EDwQPIcFLitdh33Ehy4YK119EMQAERI5OQ8PhwjEhw4QxAjEhw4QxMQIxAcOEDw8CDxZMTABQ1xYtA4YHTkLuP/eQAsdOQwiFzkDIhc5C7j/3rIhORC4/8BAChU5ASIhOQlAHDkrKysrKysrK1ldcQArXSsrAV1ZMwEBMxcWFzY3NzMBASMDJwEPAYT+meGjLhwsJbPX/pEBi93aOv7pAigB/vlHMEIz+/4M/c4BSln+XQABACH+UQPuBCYAGgH3sQICQ1RYQB0KFA8DCwMcGQ8SBgsGE0ASDyALQAwgDxgPDwJVDxkvKxrdGhjNGhkQ3RoYzQA/Pz/tEhc5MTAbsw8cAQ+4/95AbRw5KBRWD68KA0ANQA8CDyAoMDQQICgwNAcMCRIWDRgSJwsnDCcNNgw2DTUOmRELKBIoE0gWWRJZE1kVaRJpE2kVeQZ2DXkRehR6FYUNihGMEowTiRSYCqgLvBC7EboU6grnFPUN/RD5FP8cHhKxBgJDVFhAFhMLHBsED0QPhA8DDxkLAxwZDxIGCwYAPz8/7RESOV0BERI5ORtANw8PDBAREhIKAAMZFBMTJRIKFBISCg8MDxEMJQsKFAsLChMSEgwMCwYDHBkPABwQHAIvHL8cAhy4Aj+1DxNAEkAUuAJUQAs/EkASAl8SvxICErgBQrYPASIARRsKuAJUQBIPIAtAQCAMMAxPDANQDP8MAgy4AUKzLw8BD7gCP7QbIHxmGCsaGRD9cfRdcRoY7RoZEO0YEPTkGRDkXXHtGhgQ7RkQ5F1xABg/7T88EDwQPIcFLisIfRDEhwUuGCsOfRDEABESOYcOEDw8CMRLsA5TS7AYUVpYuwAM/+gAC//oATg4WVkxMAFDXFi5ABT/3rY3OQoiNzkOuP/otRU5ESIVOSsrKytZXXErKwBxXSsBXVkTJxYzMjY3Njc2NwEzExYXNjcTMwEGBwYGIyJ/FDssPEgXESYFC/5twt0rIh8r47T+bEEkMHxWNP5nqRAoJBtrDx0EKP2ZdYF8dgJr+8ivQllTAAABACgAAAPUBCYADgGvQA0SuALJCAISATISFzQIuP/OQAkSFzQBPh4hNAi4/8JASh4hNCkCKAkvEDkBOQpJAUYCRghJCU8QXAFUAlQIWglQEGwBYwJjCGoJewF0CHsJiwGFCIkJ+QH0AhsZCCYBKQgrCTkIpQjXAQcQuP/AtxAVNAIsEjkJuP/UQCMSOQECOgkKAggKCiUBAhQBAQIBDQ4IBgJhBSsHBgYKYQ0ADbj/9EAJCwsGVQ0rDgoCuAEPtAgIBwUGuwJbAAAAB//0QBYLCwZVByINoA4BAA5ADmAOgA7wDgUOuP/0QCQLCwZVDnQACn4BAa8AAU8AbwD/AAMAGAsLBlUAGQ8QdCF8xBgrK070K11xPE0Q7RD9K11xPOQrEPQ8EDwQ/QA/7Ss8EOU/PP3lETkREjmHBS4rh33EEA7EKzEwASsrK3FdACsrKytDXFi1KQEmCAIBuP/OQAkSFzQIMhIXNAG4/8K3HiE0CD4eITQAKysrKwFxWQFdQ1xYuQAI/96yDzkJuP/esg85Cbj/6LcbOQkIFhs9Cbj/8LIXOQm4//hAChY5AhQWOQIaFjkrKysrKysrK1kzNQEGIyE1IRUBBzYzIRUoAqRzWP5PA2T9wW95agHrkgMIBpJ3/V57CZsAAAMAA//uBegF0wAPAB8AOgEzQCCUEpQWmxqbHqYDqAuoDbkw1BLUFtsa2x7VM9Y2DnAIILgCq7MhhyQvuAKrszAuAS67AmAAKwA4AmJAEE8kAQ8kbyR/JO8kBCSUCDK4AmJACwArjyv/KwMrlAAYuAJisggLELgCYrIAAy+4AmKyLtMguAJisyGIBDW9AmIAJwJkAAwAHAJiswQaPBS4AmK1DBk7s3oYK04Q9E3tThD2Te0Q9O0Q9O307QA/7T/tEPRd7RD0XXHtEP1d5BD95DEwQ3lAVDM3JSoBHykmEiUOJgIlHiYWJgolBiYaJTMqNR8ANyU1HwARDxQhAB8BHCEBFwkUIQAZBxwhATQoMh8BNiY4HwATDRAhAR0DECEBFQsYIQAbBRghACsrKysrKwErKysrKysrKysrKysrKyuBgYEBXQEyBBIVFAIEIyIkAjU0EiQXIgQCFRQSBDMyJBI1NAIkExcGBiMiJjU0NjYzMhYXByYmIyIGFRQWMzI2Ava+AWrKx/6ZxMT+mcjLAWq+n/7TqqcBLKOjASymqf7SVHsew4uw3GS5d4WwIHcedU9zlY1wWogF08P+lcXD/pjHxwFow8UBa8N9o/7RpKP+1aenASujpAEvo/0QJH2V5MqEw2N/bR1KT6SZmZ1oAAABAGwD6QE9BckACwB0QCbTB+MHArEHwwcC8ggBkwihCAJzCIIIAlUIZQgCAggBCAsDAAirB7gBUEAeAQP5AgIBCwA8AQACAzwABzgIJwAAIAEBARkMnXkYK04Q9F08TRD05BD9PAA//TwQPBDtEP3tARESOQDJMTAAcnFxcXEBcXETNTMVFAcGByc2Njd8wR8rWyw2NQME+NGlhjtRKUcWX1MAAAAAAQAAAAU1wwAAAABfDzz1CDsIAAAAAACi4ycqAAAAANH4y3f6r/1nEAAIDAAAAAkAAQABAAAAAAABAAAHPv5OAEMQAPqv+noQAAABAAAAAAAAAAAAAAAAAAANXQYAAQAAAAAAAjkAAAI5AAACOQCwAtcAXgRzABUEcwBJBx0AdwVWAFgBhwBaAqoAfAKqAHwDHQBABKwAcgI5AKoCqgBBAjkAugI5AAAEcwBVBHMA3wRzADwEcwBWBHMAGgRzAFUEcwBNBHMAYQRzAFMEcwBVAjkAuQI5AKoErABwBKwAcgSsAHAEcwBaCB8AbwVW//0FVgCWBccAZgXHAJ4FVgCiBOMAqAY5AG0FxwCkAjkAvwQAADcFVgCWBHMAlgaqAJgFxwCcBjkAYwVWAJ4GOQBYBccAoQVWAFwE4wAwBccAoQVWAAkHjQAZBVYACQVWAAYE4wApAjkAiwI5AAACOQAnA8EANgRz/+ECqgBZBHMASgRzAIYEAABQBHMARgRzAEsCOQATBHMAQgRzAIcBxwCIAcf/ogQAAIgBxwCDBqoAhwRzAIcEcwBEBHMAhwRzAEgCqgCFBAAAPwI5ACQEcwCDBAAAGgXHAAYEAAAPBAAAIQQAACgCrAA5AhQAvAKsAC8ErABXBVb//QVW//0FxwBoBVYAogXHAJwGOQBjBccAoQRzAEoEcwBKBHMASgRzAEoEcwBKBHMASgQAAFAEcwBLBHMASwRzAEsEcwBLAjkAvQI5ACMCOf/lAjkACQRzAIcEcwBEBHMARARzAEQEcwBEBHMARARzAIMEcwCDBHMAgwRzAIMEcwBJAzMAgARzAGsEcwAbBHMAUQLNAG0ETAABBOMAmQXlAAMF5QADCAAA4QKqAN4CqgA9BGQATggAAAEGOQBTBbQAmgRkAE4EZABNBGQATQRz//0EnACgA/QAOAW0AHoGlgChBGQAAAIxAAAC9gAvAuwALQYlAH8HHQBEBOMAgQTjAJ4CqgDoBKwAcgRkAFQEcwAuBGQAMwTlABoEcwCGBHMAjAgAAO8FVv/9BVb//QY5AGMIAACBB40AUgRz//wIAAAAAqoAUwKqAEcBxwCAAccAbARkAE4D9AAvBAAAIQVWAAYBVv45BHP/5AKqAFwCqgBcBAAAFwQAABcEcwBJAjkAuQHHAGwCqgBHCAAAJQVW//0FVgCiBVb//QVWAKIFVgCiAjkAjQI5/+ACOQAEAjkAFQY5AGMGOQBjBjkAYwXHAKEFxwChBccAoQI5AMYCqgAZAqoABgKqAB0CqgAuAqoA5QKqAKICqgBrAqoAOgKqAEsCqgAoBHMAAAHHAAMFVgBcBAAAPwTjACkEAAAoAhQAvAXH//0EcwBJBVYABgQAACEFVgCeBHMAhwSsAHIErAChAqoAawKqABkCqgAhBqwAawasAGsGrAAhBHMAAAY5AG0EcwBCAjkAsQVWAFwEAAA/BccAZgQAAFAFxwBmBAAAUARzAEYEa//hAqoA7gVW//0EcwBKBVb//QRzAEoFxwCeBOsARwXH//0FVgCiBHMASwVWAKIEcwBLBHMAlgHHAEIEcwCWAlUAiARzAJoCrACDBccAnARzAIcFxwCcBHMAhwY5AGMEcwBEBccAoQKqAIUFxwChAqoAPAVWAFwEAAA/BOMAMAI5ACQE4wAwAwAAIwXHAKEEcwCDBccAoQRzAIME4wApBAAAKATjACkEAAAoBGgApAY5AGAGYgBVBKAASAR0AEgDkQBiBPAARAMpAC4FMABIBGv/4QQAALAC6wBSCMAAMwgAAE8EAACZCAAATwQAAJkIAABPBAAAmAQAAJgH1QFqBcAAngSrAHIE1QCdBKwAcQTVAiIE1QEFBav/6QUAAckFqwJ+Bav/6QWrAn4Fq//pBasCfgWr/+kFq//pBav/6QWr/+kFq//pBasBwAWrAn4FqwHABasBwAWr/+kFq//pBav/6QWrAn4FqwHABasBwAWr/+kFq//pBav/6QWrAn4FqwHABasBwAWr/+kFq//pBav/6QWr/+kFq//pBav/6QWr/+kFq//pBav/6QWr/+kFq//pBav/6QWr/+kFq//pBav/6QWr/+kFqwLWBasAZgWr/+oF1f//BNUAkggAAAAH6wEwB+sBIAfrATAH6wEgBNUAsgTVAIAE1QAqCCsBmAhrAbgHVQAQBgAA9AYAAG8EQAA6BUAANwTAAD8EFQBABAAAJQYAAFUF4QC/A40AiQTV/9kBgACAAtUAhgcVAGEClgAPBNUAkgLWAIMC1gCDBNUAsgLWAHAFVv/9BHMASgXHAGYEAABQBccAZgQAAFAFVgCiBHMASwVWAKIEcwBLBVYAogRzAEsGOQBtBHMAQgY5AG0EcwBCBjkAbQRzAEIFxwCkBHMAhwXHAB8EcwAGAjn/zgI5/84COf/kAjn/5AI5//YCOf/1AjkASwHHABkEAAA3Acf/ogVWAJYEAACIBAAAhgRzAJYBx//6BccAnARzAIcFyQClBHMAiwY5AGMEcwBEBjkAYwRzAEQFxwChAqoAawVWAFwEAAA/BOMAMAI5AAwFxwChBHMAgwXHAKEEcwCDBccAoQRzAIMFxwChBHMAgweNABkFxwAGBVYABgQAACEBxwCJBVb//QRzAEoIAAABBx0ARAY5AFME4wCBAjkAuQeNABkFxwAGB40AGQXHAAYHjQAZBccABgVWAAYEAAAhAccAigKq/+EEcwAbBM0AWgasAGsGrAAiBqwAIgasAEoCqgDiAqoAawKqAN4Cqv/qBVf//wZG/6cGtP+oAxL/qAYy/6cG2P+nBgX/pwHH/3gFVv/9BVYAlgVY//4FVgCiBOMAKQXHAKQCOQC/BVYAlgVYAAsGqgCYBccAnAUzAG0GOQBjBccApAVWAJ4E8gCUBOMAMAVWAAYFVgAJBq8AfwX7AGECOQAEBVYABgSgAEgDkQBiBHMAiwHHAGsEYACIBJoAjAQAABkDhwBIBHMAiwRzAFwBxwCJBAAAhgQAABgEnACgBAAAGgOVAFwEcwBEBI0AgwPbAFYEYACIBDMAEQW0AHoGPwBXAcf/yQRgAIgEcwBIBGAAiAY/AFcFVwCiBusAMgRVAKEFwABkBVYAXAI5AL8COQAEBAAANwh1AA0IFQCkBtUAMQSpAKEFFQAKBcAAoAVW//0FQACnBVYAlgRVAKEFawAABVYAogdjAAcE1QBOBcAAoQXAAKEEqQChBUAAEgaqAJgFxwCkBjkAYwXAAKAFVgCeBccAZgTjADAFFQAKBhUAUgVWAAkF6wCfBVUAVwdVAKEHgAChBlUAAAcVAKgFQAClBcAAVQgVAKQFxwAaBHMASgSVAFsEQACIAusAiASrAAAEcwBLBVr/+wOrADIEeACHBHgAhwOAAIYEqwAYBYAAjARrAIgEcwBEBFUAiARzAIcEAABQA6oAJgQAACEGlQBLBAAADwSVAIoEKwBFBmsAjQaVAI0FAAAoBcAAiwQrAIQEFQAwBgAAiQRVAB8EcwBLBHMAAALrAIkEFQBLBAAAPwHHAIgCOQAJAcf/ogdAABMGgACDBHMAAAOAAIYEAAAhBGsAiAPpAKEDSgCICAAAQQiVAKAFhQAtAAABAQAAAB4AAAAxAAAAMQAAAQEAAAB+AAAAfgAAAIwAAACMAAABAQAAABAAAAEBAAABIQMQAH0AAACMAjMA0gAAAwsAAP8EAjkAuQSBAGkEVgAyAzEAGQQRAC0E0QCWAfkAmwMPAF8EygCbBLgAjAH5AJsEEwAoA7AAUAO0ADwEygCbBM8AUAH5AJsC0gA8BJgAWgQ8ABkEiABuBF8AcwOxABkD1AAKBGYAlgQTACgFjgBkBSQAKAPyAJsD8gCbA/IAmwHjAFoDVgBaBoYAmwH5/6wEEwAoBBMAKAO0/1cDtP9XBEgALQWOAGQFjgBkBY4AZAWOAGQEgQBpBIEAaQSBAGkEVgAyAzEAGQQRAC0E0QCWAksAAANKAAAEuACMAksAAAQTACgDsABQA7QAPATPAFAC0gA8BJgAWgSIAG4EXwBzA9QACgRmAJYEEwAoBY4AZAUkACgB+QCbBFYAMgOwAFAEXwBzBJsAPAAA/9wAAP8lAAD/3AAA/lECjQCrAo0AoALaAEMDTQB5Aaj/ugAAAEYAAABGAAAARgAAAEYAAABIAAAARgAAAEYAAABGBDUBfAQ1AS4ENQC3BDUAgQQ1ASwENQC+BDUArwQ1AIEENQCaBDUA2wQ1AIUCjQDBBDUAswYAAQAGAAEAAkIANgYAAQAENQCeBDUAmAQ1AMsGAAEABgABAAYAAQAGAAEABgABAAAAAEYGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAUb/7oGAAEABgABAAYAAQAFtQA6BbUAOgH0/7oB9P+6BgABAAYAAQAGAAEABgABAASBADYENQA2BD3/ugQ9/7oD6QBKA+kASgZ/ABQHdgAUAyf/ugQe/7oGfwAUB3YAFAMn/7oEHv+6BRsAMgS1ACQDAP/3BgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEAAAAAMAAAAEYAAABGAAAAQAAAAEYGAAEABgABAAAA/9wAAP5RAAD/FgAA/xYAAP8WAAD/FgAA/xYAAP8WAAD/FgAA/xYAAP8WAAD/3AAA/xYAAP/cAAD/IAAA/9wEcwBKCAAAAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQACjQB/Ao0AXQYAAQAE7gAVA00AeQGoAA4B1v/cAagAVgHWABADdQAyA3UAMgGoAC0B1gATBRsAMgS1ACQB9P+6AfT/ugGoAJMB1gATBbUAOgW1ADoB9P+6AfT/ugJCAAADAP/3BbUAOgW1ADoB9P+6AfT/ugW1ADoFtQA6AfT/ugH0/7oEgQA2BDUANgQ9/7oEPf+6BIEANgQ1ADYEPf+6BD3/ugSBADYENQA2BD3/ugQ9/7oCswBfArMAXwKzAF8CswBfA+kASgPpAEoD6QBKA+kASgaSAD4GkgA+BD//ugQ//7oGkgA+BpIAPgQ//7oEP/+6CMkAPgjJAD4Gxf+6BsX/ugjJAD4IyQA+BsX/ugbF/7oEp/+6BKf/ugSn/7oEp/+6BKf/ugSn/7oEp/+6BKf/ugRaACoDmgA2BDX/ugMn/7oEWgAqA5oANgQ1/7oDJ/+6Bk8AJwZPACcCJP+6Ahr/ugSnAEYEpwBGAiT/ugIa/7oEzwAtBM8ALQMn/7oDJ/+6BA0ARwQNAEcBqP+6Aaj/ugK0ACMCtAAjAyf/ugMn/7oENQBFBDUARQH0/7oB9P+6AkIANgMA//cDmv+6Ayf/ugN1ADIDdQAyBRsAMgS1ACQFGwAyBLUAJAH0/7oB9P+6BFoAQATOAEkEWgAmBM4AOQRaAFMEzgBKBFoAUwTOAEoGAAEABgABAAAAAEYAAABGBgABAAYAAQAGAAEAAAAARgAAAEYGAAEABgABAAAAAEgAAABGBgABAAYAAQAGAAEAAAAARgAAAEYAAABGAAAARgAAAEAAAAAwBgABAAAAAEYAAABGBgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEAAo0AygKNAMcCjQDGBgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEABgABAAYAAQAGAAEAAQD/uggA/7oQAP+6BtwAYwU/AEQG1QChBVsAgwAA/dwAAPwvAAD8pgAA/lQAAPzXAAD9cwAA/ikAAP4NAAD9EQAA/GcAAP2dAAD79QAA/HIAAP7VAAD+1QAA/wIEGwCgBqwAawasABkAAP62AAD9cwAA/ggAAPymAAD+UwAA/REAAPvIAAD69AAA+q8AAPxyAAD7qgAA+2oAAPzxAAD8fQAA+90AAPzBAAD7mAAA/eoAAP6EAAD9wgAA/PEAAP1fAAD+dgAA/rwAAPzrAAD9bAAA/VgAAPyQAAD9FQAA/CwAAPwTAAD8EgAA+5YAAPuWAccAiAVW//0EcwBKBVb//QRzAEoFVv/9BHMASgVW//0EcwBKBVb//QRzAEoFVv/9BHMASgVW//0EcwBKBVb//QRzAEoFVv/9BHMASgVW//0EcwBKBVb//QRzAEoFVv/9BHMASgVWAKIEcwBLBVYAogRzAEsFVgCiBHMASwVWAKIEcwBLBVYAogRzAEsFVgCiBHMASwVWAKIEcwBLBVYAogRzAEsCOQBjAccAHwI5ALoBxwB8BjkAYwRzAEQGOQBjBHMARAY5AGMEcwBEBjkAYwRzAEQGOQBjBHMARAY5AGMEcwBEBjkAYwRzAEQG3ABjBT8ARAbcAGMFPwBEBtwAYwU/AEQG3ABjBT8ARAbcAGMFPwBEBccAoQRzAIMFxwChBHMAgwbVAKEFWwCDBtUAoQVbAIMG1QChBVsAgwbVAKEFWwCDBtUAoQVbAIMFVgAGBAAAIQVWAAYEAAAhBVYABgQAACEFVv/9BHMASgI5/+IBx/+wBjkAYwRzAEQFxwChBHMAgwXHAKEEcwCDBccAoQRzAIMFxwChBHMAgwXHAKEEcwCDAAD+/gAA/v4AAP7+AAD+/gRV//0C6wAMB2MABwVa//sEqQChA4AAhgSpAKEDgACGBccApARrAIgEc//9BAAAFARz//0EAAAUBVYACQQAAA8FVQBXBCsARQVVAKEEcwCHBgUAYwRzAFUGOQBgBHMARAW1ADoB9P+6AiT/ugIa/7oEpwBGAfQAngH0ABAB9AAbAfQAEAH0AGsB9P/5Aif/zgAAAA8AAP/1AqoApAKqAKQAAAAOAAAAVgAAAFYAAP/PAagADwHW/78BqP/1Adb/zQGoAB0B1v/1AagAkwHWABMDdQAyA3UAMgN1ADIDdQAyBRsAMgS1ACQFtQA6BbUAOgH0/7oB9P+6BbUAOgW1ADoB9P+6AfT/ugW1ADoFtQA6AfT/ugH0/7oFtQA6BbUAOgH0/7oB9P+6BbUAOgW1ADoB9P+6AfT/ugW1ADoFtQA6AfT/ugH0/7oFtQA6BbUAOgH0/7oB9P+6BIEANgQ1ADYEPf+6BD3/ugSBADYENQA2BD3/ugQ9/7oEgQA2BDUANgQ9/7oEPf+6BIEANgQ1ADYEPf+6BD3/ugSBADYENQA2BD3/ugQ9/7oEgQA2BDUANgQ9/7oEPf+6ArMAMgKzADICswBfArMAXwKzAF8CswBfArMAMgKzADICswBfArMAXwKzAF8CswBfArMAXwKzAF8CswA4ArMAOAKzAEkCswBJA+kASgPpAEoD6QBKA+kASgPpAEoD6QBKA+kASgPpAEoD6QBKA+kASgPpAEoD6QBKA+kASgPpAEoD6QBKA+kASgaSAD4GkgA+BD//ugQ//7oGkgA+BpIAPgQ//7oEP/+6BpIAPgaSAD4EP/+6BD//ugjJAD4IyQA+BsX/ugbF/7oIyQA+CMkAPgbF/7oGxf+6BKf/ugSn/7oEWgAqA5oANgQ1/7oDJ/+6Bk8AJwZPACcGTwAnAiT/ugIa/7oGTwAnBk8AJwIk/7oCGv+6Bk8AJwZPACcCJP+6Ahr/ugZPACcGTwAnAiT/ugIa/7oGTwAnBk8AJwIk/7oCGv+6BKcARgSnAEYEpwBGBKcARgk+ADIJPgAyB0D/ugdA/7oGfwAUB3YAFAMn/7oEHv+6BM8ALQTPAC0DJ/+6Ayf/ugTPAC0EzwAtAyf/ugMn/7oEzwAtBM8ALQMn/7oDJ/+6Bn8AFAd2ABQDJ/+6BB7/ugZ/ABQHdgAUAyf/ugQe/7oGfwAUB3YAFAMn/7oEHv+6Bn8AFAd2ABQDJ/+6BB7/ugZ/ABQHdgAUAyf/ugQe/7oEDQBHBA0ARwGo/7oBqP+6BA0ARwQNAEcBqP+6Aaj/ugQNAEcEDQBHAaj/ugGo/7oEDQBHBA0ARwGo/7oBqP+6BDUARQQ1AEUB9P+6AfT/ugQ1AEUENQBFBDUARQQ1AEUENQBFBDUARQH0/7oB9P+6BDUARQQ1AEUEgQA2BDUANgQ9/7oEPf+6AkIANgMA//cDGgAaAxoAGgMaABoDdQAyA3UAMgN1ADIDdQAyA3UAMgN1ADIDdQAyA3UAMgN1ADIDdQAyA3UAMgN1ADIDdQAyA3UAMgN1ADIDdQAyBRv/ugS1/7oFGwAyBLUAJAH0/7oB9P+6A3UAMgN1ADIFGwAyBLUAJAH0/7oB9P+6BRsAMgS1ACQGfwBFBn8ARQZ/AEUGfwBFAagAKAAA/ikAAP6iAAD/MAAA/x0AAP8SAAD/kgAA/n4I/AAyCK0AMgAA/7UAAP+2AAD+7QAA/2QAAP5+AAD/nwGNAAAC9v/9AAD+ggAA/xAEzQAyAAD/WAAA/1gAAP9kBpIAPgaSAD4EP/+6BD//ugjJAD4IyQA+BsX/ugbF/7oEWgAqA5oANgQ1/7oDJ/+6A00AeQK0ACMCQgA2AfT/ugKQ/7oB9AAvAfQAOwH0ABIB9ACxAfQAbQZ/ABQHdgAUAfkAmwAA/tkCvAAAA/IAmwRa//UEzv/1BFoAUwTOAEoEWgBTBM4ASgRaAFMEzgBKBFoAUwTOAEoEWgBTBM4ASgRaAFMEzgBKBDUAcQQ1AK0EWgAPBM4ADwRzABQGEQAUBUAApwRzAIYFQAAKBHMACgXHAFEFxwBmBAAAUAXH//0GegAUBUAASgRzAEYEdABIBVYAbgTVAFME4//EBjkAbQT+AA8HDACHAccAgwI5AB8FVgCWBAAAiAHHABUEAAAYByAApAXH/7gEcwCLBjkAYAbyAGMFVwBEBgkAFARzAIYFVgCeBVYAawQAAE8E8gCUAwsARAI5ACQE4wAUAjkAJATjADAF+wBhBccAoQYuABAEAAAhBOMAKQQAACgE4wApBOMAMQRcAEQEXAA/BHMAPARzAFUDqwAyA+UAJARzAIcCFAC8A04AvASsAHICOQCwCqoAngnHAJ4IZABGCH8AlgaqAJYDnACDCccAnAeOAJwGKwCHBHMAVQVW//0EcwBKAAD+/gVW//0EcwBKCAAAAQcdAEQGOQBtBHMAGgY5AG0EcwBCBVYAlgQAAIgGOQBjBHMARAY5AGMEcwBEBOMAKQRcAEwBx/+iCqoAngnHAJ4IZABGBjkAbQRzAEIIRgCkBPIAngXHAJwEcwCHBVb//QRzAEoFVv/9BHMASgVWAKIEcwBLBVYAogRzAEsCOf+KAjn/ZAI5AAQCOf/2BjkAYwRzAEQGOQBjBHMARAXHAKECqv/MBccAoQKqAGgFxwChBHMAdgXHAKEEcwCDBVYAXAQAAD8E4wAwAjkAJARcAFEDfgATBccApARzAIcFpgCkBNYAXgSGAF4E4wApBAAAKAVW//0EcwBKBVYAogRzAEsGOQBjBHMARAAA/v0GOQBjBHMARAY5AGMEcwBEBjkAYwRzAEQFVgAGBAAAIQRzAFcEcwBIBHMAhgRzAIYEAAATBAAAUARzAEYEcwBGBHMAVQXpAFUDqwBJA6sAMgUNADIEDwBEAjn/uQRzAEIEcwBCBHgAUAQCABkE7wAZBHMAiwRzAIcEcwCHAccAGQHHAFcC2QBEAp4AAAJuABQBxwCDBJMAgwaqAIQGqgCEBqoAhwRz/6YEcwCLBGwAhwRzAEQGUwBEBj8AVwRmAEQCqv/kAqr/5AKq/+QCqgCFAqoAhQKqAIUCqv/kBFUAigRVAIoEAAA/Acf/ogIU/7kBx/9yAssAAAI5AA8COQAkBHMAGQSMAFQEYACIBAAAGgXHAAYEAAAYBCgAGQQAACgEVAAoBFwATARcAHkEAAAkBAAAUAQAACQEAABQBjkAYwRAAIgEDwBJBHgAUARrAIgDLgAABAAACAM7AIgEcwBIBAAAJAQAAFAHtwBGB0AARggLAEYFswAkA28AJAXAACQGHAATBUoAgwUPAIMD4gAeBDgAYwMRAGQDEQBkAUb/zgHrAGQB6wAAAesAAALqAGQD2QAAApEAAAGHAFoC1wBeAccAgAHHAGwBxwCKAqoA+wKqAPsCygAyAsoAMgSsAHAErABwBKwAZQSsAGUCqgEhAqoA3gKqAFkCqgEhAqoAHQKqAFkCqgDeAjkAtgI5ALYCqgD7AqoA+wKqAKYCqgCmAqoApgKqAB0Cqv/iAqr/+wKUAAABQgBkArgAMgKgAAACygAyAxAAlgMQAJYDEACWAxAAlgMQAJYCqgBiAqoAYgKqACgCqgAdAqoARwRXAJYEVwCWBFcAlgRXAJYEVwBDBFcAQwRXAEMEVwBDBFcAQwMQAEMEVwAvBFcALwRXAC8EVwAvBFcALwMQAC8EVwAlBFcAJQRXACUEVwAlBFcAJQMQAC8EVwAaBFcAGgRXABoEVwAaBFcAGgMQABoEVwBCBFcAQgRXAEIEVwBCBFcAQgMQAEIEVwCWBFcAlgRXAJYEVwCWBFcAQgRXAEIEVwBCBFcAQgRXAEIDEABCBFcALwRXAC8EVwAvBFcALwRXAC8DEAAvBFcALwRXAC8EVwAvBFcALwRXAC8DEAAvBFcAJgRXACYEVwAmBFcAJgRXACYDEAAmBFcAQgRXAEIEVwBCBFcAQgRXAEIDEABCBFcAlgRXAJYEVwCWBFcAlgRXAEIEVwBCBFcAQgRXAEIEVwBCAxAAQgRXACYEVwAmBFcAJgRXACYEVwAmAxAAJgRXACMEVwAjBFcAIwRXACMEVwAjAxAAIwRXAC8EVwAvBFcALwRXAC8EVwAvAxAALwRXAEsEVwBLBFcASwRXAEsEVwBLAxAASwRXAJYEVwCWBFcAlgRXAJYEVwBCBFcAQgRXAEIEVwBCBFcAQgMQAEIEVwAaBFcAGgRXABoEVwAaBFcAGgMQABoEVwAkBFcAJARXACQEVwAkBFcAJAMQACQEVwAvBFcALwRXAC8EVwAvBFcALwMQAC8EVwBOBFcATgRXAE4EVwBOBFcATgMQAE4EVwCWBFcAlgRXAJYEVwCWAAD+wQAA/sYAAP2sAAD+2AAA/5IAAP7pAAD/TAAA/qAAAP7EAAD/zgAA/2YAAP6gAAD+2AAA/tgAAP+XAAD/mAAA/5kAAP/0AAD/QgAA/0IAAP9EAAD/XwAA/ocAAP/sAAD/pgAA/1EAAP9RAAD/UQAA/skAAP8cAAAAAAAA/ukAAP9MAAD/kwAA/yoAAP9WAAD/zgAA/ocAAP67AAD+xAAA/sQAAP7YAAD+2AAA/rMAAP7JAAD9rQAA/sgAAP6zAAD+yQAA/a0AAP4WAAD+5gAA/6YAAP6HAAD/RAAA/roAAP8jAAD/mgAA/awAAP6IAAAAAAAA/rAAAP+YAAD+kwAA/6YAAP6HAAD+HAAA/2YAAP9EAAD+sAAA/rAAAP6wAAD/AwAA/1IAAP0fAAD/UwAA/1MAAP9TAAD+tQAA/rUAAP/DAAD+rgAA/twAAP7HAAD+yAAA/twAAP4eAAD/QgAA/1EAAP63AAD+sAKqAN4CqgBZAqoA+gSaAHAEYAAABi4AFAeqAAAGLgAUBHsATAY/AFcEzwBEBjkAYwRzAEQFxwBwBAAAUATjAKgDOwCIBP8AAAQ8ADIGDQAKBJ0AQgcgAKQGqgCEBWUAYwRzAIsFZACkBAAACgVWAGsFVgBrBOAABQTFABkF5QBfBG4ARAO2ABQDRwAoBM8ARASVAFsEAABQAcf/ogY5AGADiQBNA4kAUAVWAKIFwAChBHMASwR4AIcKtABtBP4AEAY5ABQE5wAUB5kAvwW1AIgFWAABBAAABgcuAL8FkACIBqEAeAV7AHoIbQC/BvAAiATVAGYDqwAfBl8AOQWCAEgGOQBgBHMARAZtAAkFDAAaBm0ACQUMABoImABjBywARAaqACAE5gAcCYcAbQbQAFAAAP43CrQAbQT+ABAFxwBmBAAAUAQHABQAAP6mAAD+vAAA/5gAAP+YAAD8KwAA/EwFwAChBHgAhwVAAAQEKwAUBVYAngRzAIcFXQCkBGQAiATVAE4DqwAyBKkABAOAAAAF7wApBEkAKAcJAKQFLwCICRgAoAb2AIgGBgA+BCsAIwXHAGYEAABQBOMAMAOqACYHZwAxBYcAJgVVAFcEKwBFBuQACgVUAAoG5AAKBVQACgI5AL8HYwAHBVr/+wVXAKEEaACGBUAAEgSrABgFxwCkBGsAiAXHAKQEawCIBVUAVwQrAEUGqgCYBYAAjAKqAC4FVv/9BHMASgVW//0EcwBKCAAAAQcdAEQFVgCiBHMASwYFAGMEcwBVB2MABwVa//sE1QBOA6sAMgTVAE4EXABMBcAAoQR4AIcFwAChBHgAhwY5AGMEcwBEBjkAYARzAEQFwABKBBUAKwUVAAoEAAAhBRUACgQAACEFFQAKBAAAIQVVAFcEKwBFBxUAqAXAAIsFQABKBHMARge/AEoHAwBGB6YAZgaGAFMFTQBmBBMAUwfDABIHRwAYCEYApAcHAIgGOQBtBHgAUAX5ADAFUwAmAAD/QwAA/skAAP93AAD/sAAA/0cAAP9WAAD/dAAA/tcAAP6sAAAAAAAA/1IAAP9WAAAAAAAA/qwAAP2aAAAAAAAA/2oAAP98AAD/aQAA/1YAAP6sAAD/fwAA/1YAAP3vAAD/QwAA/2kAAP98AAAAAAAA/a4AAP+MAAABAgAA/v4AAP7+AAD+3wAA/t8AAP9YAAD/IAAA/v4FVv/9BHMASgVWAJYEcwCGBVYAlgRzAIYFVgCWBHMAhgXHAGYEAABQBccAngRzAEYFxwCeBHMARgXHAJ4EcwBGBccAngRzAEYFxwCeBHMARgVWAKIEcwBLBVYAogRzAEsFVgCiBHMASwVWAKIEcwBLBVYAogRzAEsE4wCoAjkAEwY5AG0EcwBCBccApARzAIcFxwCkBHMAhwXHAKQEcwCHBccAkwRzAGgFxwCkBHMAhwI5/98Bx/+SAjkAIAI5AAYFVgCWBAAAiAVWAJYEAACIBVYAlgQAAIgEcwCWAccAfgRzAJYBx/+5BHMAlgHH/6UEcwCWAcf/owaqAJgGqgCHBqoAmAaqAIcGqgCYBqoAhwXHAJwEcwCHBccAnARzAIcFxwCcBHMAhwXHAJwEcwCHBjkAYwRzAEQGOQBjBHMARAY5AGMEcwBEBjkAYwRzAEQFVgCeBHMAhwVWAJ4EcwCHBccAoQKqAIUFxwChAqoAhQXHAKECqgBeBccAoQKqACYFVgBcBAAAPwVWAFwEAAA/BVYAXAQAAD8FVgBcBAAAPwVWAFwEAAA/BOMAMAI5ACQE4wAwAjkAJATjADACOf//BOMAMAI5AA4FxwChBHMAgwXHAKEEcwCDBccAoQRzAIMFxwChBHMAgwXHAKEEcwCDBVYACQQAABoFVgAJBAAAGgeNABkFxwAGB40AGQXHAAYFVgAJBAAADwVWAAkEAAAPBVYABgQAACEE4wApBAAAKATjACkEAAAoBOMAKQQAACgEcwCHAjkAAwXHAAYEAAAhBHMASgHHAIkEoABIBKAASASgAEgEoABIBKAASASgAEgEoABIBKAASAVW//0FVv/9BoIAEwaCABMGggATBoIAEwaCAFYGggBWA5EAYgORAGIDkQBiA5EAYgORAGIDkQBiBh4AAAYeAAAHbAAAB2wAAAdsAAAHbAAABHMAiwRzAIsEcwCLBHMAiwRzAIsEcwCLBHMAiwRzAIsGjwAABo8AAAgfAAAIHwAACB8AAAgfAAAIH//zCB//8wHHAIEBxwCBAcf/mwHH/5sBx//rAcf/6wHH/6IBx/+iAwEAAAMBAAAEkQAABJEAAASRAAAEkQAABJH/8wSR//MEcwBEBHMARARzAEQEcwBEBHMARARzAEQGnQAABp0AAAgtAAAILQAAB8kAAAfJAAAEYACIBGAAiARgAIgEYACIBGAAiARgAIgEYACIBGAAiAaCAAAHrgAACBIAAAeuAAYGPwBXBj8AVwY/AFcGPwBXBj8AVwY/AFcGPwBXBj8AVwZfAAAGXwAAB+8AAAfvAAAHiwAAB4sAAAeL//8Hi///BKAASASgAEgDkQBiA5EAYgRzAIsEcwCLAcf/5gHHAGgEcwBEBHMARARgAIgEYACIBj8AVwY/AFcEoABIBKAASASgAEgEoABIBKAASASgAEgEoABIBKAASAVW//0FVv/9BoIAEwaCABMGggATBoIAEwaCAFYGggBWBHMAiwRzAIsEcwCLBHMAiwRzAIsEcwCLBHMAiwRzAIsGjwAABo8AAAgfAAAIHwAACB8AAAgfAAAIH//zCB//8wY/AFcGPwBXBj8AVwY/AFcGPwBXBj8AVwY/AFcGPwBXBl8AAAZfAAAH7wAAB+8AAAeLAAAHiwAAB4v//weL//8EoABIBKAASASgAEgEoABIBKAASASgAEgEoABIBVb//QVW//0FVv/9BVb//QVW//0CqgDlAqoA/QKqAOUCqgAGAqoABgRzAIsEcwCLBHMAiwRzAIsEcwCLBoIAAAaCAAAG8wAABvMAAAXHAKQCqgATAqoAEwKqAAYBx/+7Acf/qwHH/8oBx//KAcf/kwHH/5MCOQAaAjn/9QNlAAADZQAAAqoAEwKqABMCqgAGBGAAiARgAIgEYACIBGAAiASNAIMEjQCDBGAAiARgAIgFVgAGBVYABgbmAAAHGAAABh4AAAKq/+oCqv/qAqoAWQY/AFcGPwBXBj8AVwY/AFcGPwBXB2UAAAadAAAHJwAABl8AAAX7AGECqgDeAqoA5QRzAA0FxwBmBccAZgaqAIcFxwAkCVAAoQeNABkFVgAfBOMAMAgAACkEAAAwBMEAZgAA/1MAAP9TAAD/UwAA/1MBxwAZAcf/ogQrAAUFVgARBXQARgLL/6MFegCHAvD/yAV/AAoFfwAKAqoAhAKqAIQCqgDJAqoAyQKqAKACqgBZAqr/rwKqADoCqgAGAjkAuQKqAKkCqgCpAqoAqQKqAKkDLgAeAy4AHgKqADoAAP9zAAD/pQAA/tgAAP8jAAD/cgAA/3IAAP7nAAD/pQAA/1MAAP9TAAD/UwVWAJ4EcwCHA/gAGQX7ABkHHQBEBEAAGQQAAFAEaQCHBGkAGQPrAIcDqwAyAccAiANhAEEEAACIAzYAEAWAAIwEeACHBHMARAQAABME3gBEBN4ARATeAA0HjQBQA6gARARzAEQEcwBEBCsAhARVAB8EVQAfA6oAJgRgAIgExgBEBd4ARATGAEQEAAAaBccABgQAACgDqwAyA2sAPwTbAB8C6wCIBAAAGgRVAIgEKwCEBbQAegSrABgDoAAABU8AAANRADIDUf/RA5gAMgNIADIDSAAyA/gAMgNuADIBVgBpAoQALQNmADIC0AAyBBUAMgNxADIDbwAyBBgAMgMPADIDWQAyA5wAMgN2ADEDbwAyBPsAAAL6ADIC+gAyAwQAMgTMADIDBQBkAwUAMgL5ADIC+QAyAowAMgKMADIDBAAyAUIAZAK2AGQElQBkAw8AZAMFADIC1QAyAwUAMgMFADIDBgBkAcIAMgMPAGQDQgAyBJUAZAKSAAADIAAAAxUAZAKSAAADBgAyA4UAMgK/AAABQgBkAesAZAMPAGQCkgAAAxUAZAKSAAADCQAyA4UAMgK/AAAF7QBGCmYARgYTAEYGif+6BUH/ugHpADwEWgARAAD/DQAA/zUAAP7OAAD+twAA/skAAP/PAAD/TwAA/54AAP7KArMAXwKzAF8D6QBKA+kASgOa/7oDJ/+6A5r/ugMn/7oFrQBpBT0ALQX9AJYE3ABQBOAAPAX2AJsFPwAoBlAAKASsAHIAAP47AAD+ZgAA/mYEc//8AqoAUwLV/84BqP+6Aaj/ugGo/7oBqP+6BlgAFQnFAEcEAAAACAAAAAQAAAAIAAAAAqsAAAIAAAABVQAABHMAAAI5AAABmgAAAKsAAAAAAAAF5QADBccAZgaqAJgFgACMB0QAgwcYAEYHGABIBVb//QXHAGYEAAAUBHMACgTjADAEAABPBAAAKASlAB0AAAECAAD/QgAA/r8AAP86AAD/UwSNAAoFxwBRBccAZgXHAFEEVQChAusAiAAA/0MAAP8EAAD/rALSAJYAAP83Ahr/ugJQAB4AAP86AAD/WwAA/18AAP9+AAD/lAAA/0oAAP6cBbUAOgW1ADoB9P+WAfT/lgW1ADoFtQA6AfT/ugH0/7oFtQA6BbUAOgH0/7oB9P+6BbUAOgW1ADoB9P+6AfT/ugW1ADoFtQA6AfT/ugH0/7oFtQA6BbUAOgH0/7oB9P+6BbUAOgW1ADoB9P+6AfT/ugSBADYENQA2BD3/ugQ9/7oEgQA2BDUANgQ9/7oEPf+6ArMAMgKzADICswBfArMAXwPpAEoD6QBKBpIAPgaSAD4EP/+6BD//ugRaACoDmgA2BDX/ugMn/7oEWgAqA5oANgQ1/7oDJ/+6BFoAKgOaADYENf+6Ayf/ugZPACcGTwAnAiT/ugIa/7oGTwAnBk8AJwIk/7oCGv+6Bn8AFAd2ABQDJ/+6BB7/ugZ/ABQHdgAUAyf/ugQe/7oGfwAUB3YAFAMn/7oEHv+6ArQAIwK0ACMDJ/+6Ayf/ugK0ACMCtAAjAyf/ugMn/7oENQBFBDUARQH0/7oB9P+6BDUARQQ1AEUB9P+6AfT/ugQ1AEUENQBFAfT/ugH0/7oEDQBHBA0ARwGo/7oBqP+6A+kASgPpAEoD6QBKA+kASgaSAD4GkgA+BD//ugQ//7oEc/+TBHMARgI5/78Gqv/VBHP/twRz/5ECqv+kAqr/pAQA//8COf+5BAAAKARzAIkDCwBkBHQASAZJACQBxwAZAccAGQRzAB4EYAAeBIwACgRzAIYEcwBGAjkAEwW0AEIEAACIAcf//AaqAIcEcwCLBHMAhwKq//sEAAA/Axj/ogQAABoEAAAPBAAAKARzAEoEcwBIBHMARgRzAEsDqwBJA6sAMgU0AFUBxwCIBAAAEwHH/6IEcwCDBFwATAMEAGQC1QAyAskAMwL8ADICjAAyAdUAMgHVAAADBAAyAxEAZAFCABkBQgBkAUIAZAFCABkCKgAAAUIAZAFCAAkCMwBkBJMAZASTAGQDD//JAw8AZAMOAGQDBQAyAwAAMgK4ADIBQv/KAcIAMgMPAB0DGgAyAwYAZALUAGQCkgAAAt4AMgLeADIC3gAyAvQAMgLqADIAAP68AAD+vAAA/3MAAP6pAjkAuQL6ADIC+QAyAwUAMgKgAAAC+QAyBjkAbQVW//0EcwAPBccAZgKqAEEEoABIBKAASASgAEgEoABIBKAASASgAEgEoABIBKAASAHH/5sBx/+rAcf/mwHH/6sBx/+bAcf/uwHH/5sBx/+7BGAAiARgAIgEYACIBGAAiARgAIgEYACIBGAAiARgAIgBx/+rAcf/qwHH/7sBx/+7BGAAiARgAIgEYACIBGAAiARaAFMEzgBKA6AAEwVWABEFxwApBVgACwVWAKIEcwBLBAAAMwHH/6IF5gBjBHMASAXHAAACqgAPBVYABgQAACEEAAATBAAAUAQAABMBxwCDBFX//QLrAAEFVgAJBAAADwVWAAkEAAAPBNUAUwOrAEkFQAASBKsAGAAA/sYAAP7UAAD+xgAA/tQAAP5fAAD+XwAA/3IAAP9zAAD+5weLAAoD6wBMBAAAEwRzAAoBxwAVBHP/9AVWABEFxwChBHMAGQI5/4sFxwCkBHMAhwVWAJYEAACIBOMAKQQAACgEAAA7BJ4ApANnAIgFMABIAAD/UwAA/7wAAP7+AAD+/gAA/qQAAP6kAccAiAXJAKUFxwCcBckApQAA/s0AAP9IAAD+yQAA/s4AAP7FAAD+0AAA/tEAAP7uAAD+1gAA/twAAP3ZBjkAWARzAEgHjQAZBccABgWfAKQAAP65BdwAYwTGAAkITAAZBroABgI5ALkDgAByAYcAWgGHAFoEAACZBAAAmQI5ALACOQCwAjkAsAKqABkE4wAwBHMAUARzAA8EcwAcBlsAhwZKAEwAAAAAAAAAKgAAACoAAAAqAAAAKgAAACoAAAAqAAAAKgAAACoAAAHSAAAB0gAAAdIAAAJSAAAC+AAAAvgAAANgAAAD2AAABB4AAARaAAAEygAABoYAAAdiAAAJjAAAC2YAAAzGAAAOgAAAEFYAABECAAATlgAAFcoAABYmAAAWJgAAFiYAABaWAAAWlgAAF4gAABeIAAAZMgAAGsoAABwEAAAdTAAAHhAAAB7GAAAgVgAAIVwAACJAAAAjKAAAJV4AACXoAAApEgAAKrwAACvwAAAs9gAALuoAADFWAAA0AAAANK4AADXSAAA3RgAAOYQAADyQAAA+NgAAPjYAAD42AAA+NgAAPjYAAD42AAA+agAAPmoAAEE8AABDGgAARM4AAEaCAABIQAAASZQAAEuEAABNKAAAThwAAE80AABRzAAAUsgAAFT4AABWvgAAWIAAAFpEAABb2gAAXOAAAGCIAABhrAAAY0oAAGVoAABp0gAAa/YAAG5OAABwNgAAcDYAAHA2AABwNgAAcDYAAHA2AABwNgAAcDYAAHA2AABwNgAAcDYAAHA2AABwNgAAcDYAAHA2AABwNgAAcDYAAHA2AABwNgAAcDYAAHA2AABwNgAAcDYAAHA2AABwNgAAcDYAAHA2AABwNgAAcDYAAHA2AABwNgAAcDYAAHA2AABwNgAAcDYAAHA2AABwNgAAcDYAAHA2AABwNgAAcDYAAHA2AABwNgAAcDYAAHA2AABwNgAAciYAAHImAAByJgAAciYAAHImAAByJgAAciYAAHImAAByJgAAciYAAHImAAByJgAAciYAAHImAAByJgAAciYAAHImAAByJgAAciYAAHImAAByJgAAciYAAHImAAByJgAAciYAAHImAAByJgAAciYAAHImAAByJgAAciYAAHImAAByJgAAciYAAHImAAByJgAAciYAAHImAAByJgAAciYAAHImAAByJgAAciYAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygAAcsoAAHLKAAByygABAAANXQDyADwAnQAHAAIAEAAvAFYAAASs//8ABQACAAAAFAD2AAEAAAAAAAAAEAAAAAEAAAAAAAEADAAQAAEAAAAAAAIABwAcAAEAAAAAAAMADAAjAAEAAAAAAAQADAAvAAEAAAAAAAUADAA7AAEAAAAAAAYADABHAAEAAAAAAAcABwBTAAEAAAAAAAgABwBaAAEAAAAAAAkABwBhAAMAAQQJAAAAIABoAAMAAQQJAAEAGACIAAMAAQQJAAIADgCgAAMAAQQJAAMAGACuAAMAAQQJAAQAGADGAAMAAQQJAAUAGADeAAMAAQQJAAYAGAD2AAMAAQQJAAcADgEOAAMAAQQJAAgADgEcAAMAAQQJAAkADgEqT3JpZ2luYWwgbGljZW5jZUJFRk5HQStBcmlhbFVua25vd25CRUZOR0ErQXJpYWxCRUZOR0ErQXJpYWxWZXJzaW9uIDAuMTFCRUZOR0ErQXJpYWxVbmtub3duVW5rbm93blVua25vd24ATwByAGkAZwBpAG4AYQBsACAAbABpAGMAZQBuAGMAZQBCAEUARgBOAEcAQQArAEEAcgBpAGEAbABSAGUAZwB1AGwAYQByAEIARQBGAE4ARwBBACsAQQByAGkAYQBsAEIARQBGAE4ARwBBACsAQQByAGkAYQBsAFYAZQByAHMAaQBvAG4AIAAwAC4AMQAxAEIARQBGAE4ARwBBACsAQQByAGkAYQBsAFUAbgBrAG4AbwB3AG4AVQBuAGsAbgBvAHcAbgBVAG4AawBuAG8AdwBuAAAAAwAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAALkAVAMosyYYH9C8AykA4AMpAAIDKbIrHR+5AycDHbI7H0C4AyOzEhUyD0EtAyAAAQAvAyAAAQAgAyAAbwMgAK8DIAC/AyAABABfAx4AAQAQAx4AfwMeAIADHgCvAx4AvwMeANADHgAGAAADHgAQAx4AIAMeAG8DHgCfAx4A4AMeAAYDHQMcsiAfEEEnAxkAfwMZAAIADwMXAO8DFwD/AxcAAwAfAxcALwMXAE8DFwBfAxcAjwMXAJ8DFwAGAA8DFwBfAxcAbwMXAH8DFwC/AxcA8AMXAAYAQAMXspIzQLgDF7KLM0C4AxezamwyQLgDF7JhM0C4AxezXF0yQLgDF7NXWTJAuAMXs01RMkC4AxezREkyQLgDF7I6M0C4AxezMTQyQLgDF7MuQjJAuAMXsycsMkC4AxezEiUygLgDF7MKDTLAQRYDFgDQAxYAAgBwAxYAAQLEAA8BAQAfAKADFQCwAxUAAgMGAA8BAQAfAEADErMkJjKfvwMEAAEDAgMBAGQAH//AAwGyDREyQQoC/wLvABIAHwLuAu0AZAAf/8AC7bMOETKfQUoC4gCvAuIAvwLiAAMC4gLiAuEC4QB/AuAAAQAQAuAAPwLgAJ8C4AC/AuAAzwLgAO8C4AAGAuAC4ALfAt8C3gLeAA8C3QAvAt0APwLdAF8C3QCfAt0AvwLdAO8C3QAHAt0C3QAQAtwAAQAAAtwAAQAQAtwAPwLcAAIC3ALcABAC2wABAtsC2wAPAtoAAQLaAtr/wALTsjc5Mrn/wALTsisvMrn/wALTsh8lMrn/wALTshcbMrn/wALTshIWMrgC0rL5KR+5AyYDHLI7H0C7AyIAPgAzAyKyJTEfuAMYsjxpH7gC47MgKx+gQTAC1ACwAtQAAgAAAtQAEALUACAC1ABQAtQAYALUAHAC1AAGAGAC1gBwAtYAgALWAJAC1gCgAtYAsALWAAYAAALWABAC1gAgAsoAIALMACAC1gAwAtYAQALWAFAC1gAIAtCyICsfuALPsiZCH0EWAs4CxwAXAB8CzQLIABcAHwLMAsYAFwAfAssCxQAXAB8CyQLFAB4AHwLKAsayHh8AQQsCxgAAAscAEALGABACxwAvAsUABQLBsyQSH/9BEQK/AAEAHwK/AC8CvwA/Ar8ATwK/AF8CvwCPAr8ABgK/AiKyZB8SQQsCuwDKCAAAHwKyAOkIAAAfAqYAoggAQGofQCZDSTJAIENJMkAmOj0yQCA6PTKfIJ8mAkAmlpkyQCCWmTJAJo6SMkAgjpIyQCaEjDJAIISMMkAmeoEyQCB6gTJAJmx2MkAgbHYyQCZkajJAIGRqMkAmWl8yQCBaXzJAJk9UMkAgT1QyuAKetyQnHzdPawEgQQ8CdwAwAncAQAJ3AFACdwAEAncCdwJ3APkEAAAfApuyKiofuAKaQCspKh+AugGAvAGAUgGAogGAZQGAfgGAgQGAPAGAXgGAKwGAHAGAHgGAQAGAuwE4AAEAgAFAtAGAQAGAuwE4AAEAgAE5QBgBgMoBgK0BgHMBgCYBgCUBgCQBgCABN0C4AiGySTNAuAIhskUzQLgCIbNBQjJAuAIhsz0+Mg9BDwIhAD8CIQB/AiEAAwC/AiEAzwIhAP8CIQADAEACIbMgIjJAuAIhsxkeMkC4AiKzKj8yQLgCIbMuOjJvQUgCwwB/AsMAjwLDAN8CwwAEAC8CwwBgAsMAzwLDAAMADwLDAD8CwwBfAsMAwALDAO8CwwD/AsMABgDfAiIAAQCPAiIAAQAPAiIALwIiAD8CIgBfAiIAfwIiAO8CIgAGAL8CIQDvAiEAAgBvAiEAfwIhAK8CIQADAC8CIQA/AiEATwIhAAMCwwLDAiICIgIhAiFAHRAcECsQSAOPHAEPHgFPHv8eAjcAFhYAAAASEQgRuAENtvcN+PcNAAlBCQKOAo8AHQAfApACjwAdAB8Cj7L5HR+4AZiyJrsfQRUBlwAeBAEAHwE5ACYBJQAfATgAcwQBAB8BNQAcCAEAHwE0ABwCqwAfATKyHFYfuAEPsiYsH7oBDgAeBAG2H/kc5B/pHLgCAbYf6By7H9cguAQBsh/VHLgCq7Yf1ByJH8kvuAgBsh+8JrgBAbIfuiC4AgG2H7kcOB+tyrgEAbIfgSa4AZqyH34muAGath99HEcfaxy4BAGyH2UmuAGash9ec7gEAUAPH1ImWh9IHIkfRBxiH0BzuAgBth8/HF4fPCa4AZqyHzUcuAQBth8wHLsfKxy4BAG2HyocVh8pHLgBAbIfIx64BAGyH1U3uAFoQCwHlgdYB08HNgcyBywHIQcfBx0HGwcUCBIIEAgOCAwICggICAYIBAgCCAAIFLj/4EArAAABABQGEAAAAQAGBAAAAQAEEAAAAQAQAgAAAQACAAAAAQAAAgEIAgBKALATA0sCS1NCAUuwwGMAS2IgsPZTI7gBClFasAUjQgGwEksAS1RCsDgrS7gH/1KwNytLsAdQW1ixAQGOWbA4K7ACiLgBAFRYuAH/sQEBjoUbsBJDWLkAAQERhY0buQABASiFjVlZABgWdj8YPxI+ETlGRD4ROUZEPhE5RkQ+ETlGRD4ROUZgRD4ROUZgRCsrKysrKysrKysrGCsrKysrKysrKysrGCsdsJZLU1iwqh1ZsDJLU1iw/x1ZS7CTUyBcWLkB8gHwRUS5AfEB8EVEWVi5Az4B8kVSWLkB8gM+RFlZS7gBVlMgXFi5ACAB8UVEuQAmAfFFRFlYuQgeACBFUli5ACAIHkRZWUu4AZpTIFxYuQAlAfJFRLkAJAHyRURZWLkJCQAlRVJYuQAlCQlEWVlLuAQBUyBcWLFzJEVEsSQkRURZWLkXIABzRVJYuQBzFyBEWVlLuAQBUyBcWLHKJUVEsSUlRURZWLkWgADKRVJYuQDKFoBEWVlLsD5TIFxYsRwcRUSxHhxFRFlYuQEaABxFUli5ABwBGkRZWUuwVlMgXFixHBxFRLEvHEVEWVi5AYkAHEVSWLkAHAGJRFlZS7gDAVMgXFixHBxFRLEcHEVEWVi5DeAAHEVSWLkAHA3gRFlZKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKysrKytlQisrAbM7WWNcRWUjRWAjRWVgI0VgsIt2aBiwgGIgILFjWUVlI0UgsAMmYGJjaCCwAyZhZbBZI2VEsGMjRCCxO1xFZSNFILADJmBiY2ggsAMmYWWwXCNlRLA7I0SxAFxFVFixXEBlRLI7QDtFI2FEWbNHUDQ3RWUjRWAjRWVgI0VgsIl2aBiwgGIgILE0UEVlI0UgsAMmYGJjaCCwAyZhZbBQI2VEsDQjRCCxRzdFZSNFILADJmBiY2ggsAMmYWWwNyNlRLBHI0SxADdFVFixN0BlRLJHQEdFI2FEWQBLU0IBS1BYsQgAQllDXFixCABCWbMCCwoSQ1hgGyFZQhYQcD6wEkNYuTshGH4bugQAAagACytZsAwjQrANI0KwEkNYuS1BLUEbugQABAAACytZsA4jQrAPI0KwEkNYuRh+OyEbugGoBAAACytZsBAjQrARI0IAK3R1c3UAGEVpREVpREVpRHNzc3N0dXN0dSsrKyt0dSsrKysrc3Nzc3Nzc3Nzc3Nzc3Nzc3Nzc3Nzc3NzcysrK0WwQGFEc3QAAEuwKlNLsD9RWlixBwdFsEBgRFkAS7A6U0uwP1FaWLELC0W4/8BgRFkAS7AuU0uwOlFaWLEDA0WwQGBEWQBLsC5TS7A8UVpYsQkJRbj/wGBEWSsrKysrKysrKysrKysrKysrK3UrKysrKysrQ1xYuQCAAruzAUAeAXQAc1kDsB5LVAKwEktUWrASQ1xaWLoAnwIiAAEAc1kAK3RzASsBcysrKysrKysrc3NzcysrKysrACsrKysrKwBFaURzRWlEc0VpRHN0dUVpRHNFaURFaURFaURzdEVpREVpRHMrKysrK3MrACtzK3R1KysrKysrKysrKysrKytzdHVzK3N0dXN0dSsrK3QrKwAA); }&#xA;@font-face { font-family: &quot;g_font_8&quot;; src: url(data:font/opentype;base64,AAEAAAANAIAAAwBQT1MvMgRuLT0AAADcAAAAYGNtYXAAC+D/AAABPAAAACxjdnQgTw5I2QAAAWgAAAV0ZnBnbY+n6YkAAAbcAAAEI2dseWYF2+gZAAALAAAAAnJoZWFkuhmV8AAADXQAAAA2aGhlYQ4+B1QAAA2sAAAAJGhtdHjKwDzQAAAN0AAAAzRsb2Nhb4lwwgAAEQQAAAGcbWF4cAMrAWcAABKgAAAAIG5hbWW3Zg0jAAASwAAAAi5wb3N0AAMAAAAAFPAAAAAgcHJlcG6IrVkAABUQAAACegADAiQB9AAFAAACigK7AAAAjAKKArsAAAHfADEBAgAAAAAGAAAAAAAAAAAAAAAQAAAAAAAAAAAAAAAqMjEqAADgAODMBmn+ZQBkBmkBmwAAAAAAAAAAAAAAAAAA4AAAAwAAAAEAAwABAAAADAAEACAAAAAEAAQAAQAA4Mz//wAA4AD//yAAAAEAAAAABZEAAAXBAAAFGwBaBbMABAAA/+QAAAAAARX+6wAAAAAFwQAAAAAAAP/kAAAFpAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAP///////////////////////////////wAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAD///////8AAAAAADIAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAMgCVApkARgBHAQUAQAB3AEMAKABBACsA5gA5AIgALwAnALQAAwApAC0AegFHAAQBlABiBcAArADEApkCtgBVAFoCmQAoAEIAigCZAKEADQAqAEcAbgBwBbQANgA9AEcARwD+AYkBpAHoAkoCbgAFAA8AJAAqACoAjACYALAA2QDrATkBPQFyAZEBmAGiAfAFwAAfADYAOwBHAEcAUQB6AL8AwgDlAj4ACAAOABYAFgAmAEcAcQCzANkA7AFnAYgByAHpArYANgA8AEEATgBRAFYAWgCIAJUAnQCyAL8AwwDHAMgA1wEHASkBSwFLAXEBiQGSAhYCWQJZAloCcwK3BfAAFgAZACMAKQAqACoAMQA8AD8AUQBRAFUAWwB0AHYAeQCAAJcAowDBAMoA3ADwAQkBJwErASsBMwFUAWsBawGRAasBxgHhAiQCKgJBAm8CeAKuBhcAEQAnACsAMQA/AFUAYQBiAGgAaQBvAHMAfwB/AIEAhACGAJIAlwCaAJ0AnwCfAKsArgC9AM8A0gDdAPEA8gENASUBMwE4AVwBaAF8AYkBnAGdAaMBtgHQAdsB2wH8AgkCQwKSA6YEqAUVBZYGIga3BtIAEQAgADIAPAA8ADwAPQBHAFUAVgBXAFoAWwBcAFwAcQBzAHQAdQB2AHwAgACCAI0AngCxALIAsgCyALcAxADEANEA2QDcAN0A7wDyAPUA9gEBAQMBBgEHAQsBEAEWAScBLgEzATsBSgFOAVEBVQFbAV0BZAFpAXEBcgGQAZABlAGZAaMBpgGmAacBsQGzAbMBuQG7AcYBxwHIAdoB8gIaAh8CNQI3Aj0CSQJTAlMCYwJ3AoMChgKRApYClgKWAswC0ALRAtQC5wL8AwkDKAM2AzsDZAN0A6MDywQ3BDkEoATVBNoE3ATcBNwE6QT+BR4FOAVYBYEFlgXYBd0GEwZkBqIGtgbWBt8G6Ab6B4cADQAkAEMAVQBaAG4AcgB9AIoAiwCPAJcApgCpALYAtgC3AMQAzwDTANoA2wDlAOUA6wDuAQsBFQEcASABRgFGAUYBSQFZAVoBbQFyAXUBdgF+AZEBkgGcAaYBpwGpAcEBwwHFAd4B3wHhAfIB8wH5Af0B/QIAAhUCFgIZAhoCHgIfAiICLwI0AjQCPQJIAloCWgJdAmQCbgJ4AoECgQKIApACpgKoAqsCvwLDAsQCywLcAuAC8AL7AwsDDwMmAysDNAM1A1wDcgOLA40DngOgA6QDrQPGA9ED0QPZA/sEAARQBHoEjgTZBQAFAQUVBTYFXwWCBaIFuQXmBe8GCwYVBhoGHQYxBkkGSgZVBmsGfgaXBsgG9gcDBxYHLAdJB4cHxwCPAJ0AjQAAAAAAAAAAAAAAAAAAAHIATQCnAFwBmwAoACsAAQAiALkEWwBlAx4ChQFZAMID/ADCA/wAmwEoAH4AvQESBDcASwCpASsAfgFfAZgASgBXBcAAnQFkAMcA2gB8AD0AsgG/AB4DJgE6ANgAAgAtANkAlQEcAL8CBwKuBY4BqQCJADwA+ABHADUAbgO9A9UDuwJYAGsA8AGuAQUANwHUA1wBbgHHAwoCYgLwAtoDXAE4BP4F7wXBAAABGAA8Au0CsgC1ACACkwJeBH0DLkA1NDMyMTAvLi0sKyopKCcmJSQjIiEgHx4dHBsaGRgXFhUUExIREA8ODQwLCgkIBwYFBAMCAQAsRSNGYCCwJmCwBCYjSEgtLEUjRiNhILAmYbAEJiNISC0sRSNGYLAgYSCwRmCwBCYjSEgtLEUjRiNhsCBgILAmYbAgYbAEJiNISC0sRSNGYLBAYSCwZmCwBCYjSEgtLEUjRiNhsEBgILAmYbBAYbAEJiNISC0sARAgPAA8LSwgRSMgsM1EIyC4AVpRWCMgsI1EI1kgsO1RWCMgsE1EI1kgsAQmUVgjILANRCNZISEtLCAgRRhoRCCwAWAgRbBGdmiKRWBELSwBsQsKQyNDZQotLACxCgtDI0MLLSwAsEYjcLEBRj4BsEYjcLECRkU6sQIACA0tLEWwSiNERbBJI0QtLCBFsAMlRWFksFBRWEVEGyEhWS0ssAFDYyNisAAjQrAPKy0sIEWwAENgRC0sAbAGQ7AHQ2UKLSwgabBAYbAAiyCxLMCKjLgQAGJgKwxkI2RhXFiwA2FZLSxFsBErsEcjRLBHeuQYLSy4AaZUWLAJQ7gBAFRYuQBK/4CxSYBERFlZLSyKA0WKioewESuwRyNEsEd65BgtLC0sS1JYIUVEGyNFjCCwAyVFUlhEGyEhWVktLAEYLy0sILADJUWwSSNERbBKI0RFZSNFILADJWBqILAJI0IjaIpqYGEgsBqKsABSeSGyGkpAuf/gAEpFIIpUWCMhsD8bI1lhRByxFACKUnmzSUAgSUUgilRYIyGwPxsjWWFELSyxEBFDI0MLLSyxDg9DI0MLLSyxDA1DI0MLLSyxDA1DI0NlCy0ssQ4PQyNDZQstLLEQEUMjQ2ULLSxLUlhFRBshIVktLAEgsAMlI0mwQGCwIGMgsABSWCOwAiU4I7ACJWU4AIpjOBshISEhIVkBLSxFabAJQ2CKEDotLAGwBSUQIyCK9QCwAWAj7ewtLAGwBSUQIyCK9QCwAWEj7ewtLAGwBiUQ9QDt7C0sILABYAEQIDwAPC0sILABYQEQIDwAPC0ssCsrsCoqLSwAsAdDsAZDCy0sPrAqKi0sNS0sdrBLI3AQILBLRSCwAFBYsAFhWTovGC0sISEMZCNki7hAAGItLCGwgFFYDGQjZIu4IABiG7IAQC8rWbACYC0sIbDAUVgMZCNki7gVVWIbsgCALytZsAJgLSwMZCNki7hAAGJgIyEtLLQAAQAAABWwCCawCCawCCawCCYPEBYTRWg6sAEWLSy0AAEAAAAVsAgmsAgmsAgmsAgmDxAWE0VoZTqwARYtLEUjIEUgsQQFJYpQWCZhiosbJmCKjFlELSxGI0ZgiopGIyBGimCKYbj/gGIjIBAjirFLS4pwRWAgsABQWLABYbj/wIsbsECMWWgBOi0ssDMrsCoqLQAAAgEAAAAFAAUAAAMABwAqtQSQAAeQAbgCNLIACgS+AToAAAAFAToAAwIvAAAv/uUQ5QA//uUQ5TEwIREhESUhESEBAAQA/CADwPxABQD7ACAEwAAAAQAk/+wFxgWlAB8AKrIAAB26AgIABwI7tBMJAAAJuAI6sxoaISAREjkv7Rk5LwAYP+3tOS8xMAE2EgA+AjMyFRQGBwYAAwYHBiMiJicmJyY1NDYzMhYB32HgAQKINLIhFQ8ktf5OkjsWFnVUITJSazZ2JzKSARPaAZUBbIcXGRAKEyCo/XD+l5AdHiJMf3E5HShTbgAAAf///4kEigUbAFcAgkA0CQk+PjATFQ8PFRUGMDBCBgRCKiUoPj4ACQkAACADDxMaAxIlJSgSElkMLSAuLiggQkJUILgB8bIDAyi4AimzVFRZWBESOS/tOS/tEjkvERI5LxI5OREzLxI5LxIXORESOS8ZOS8SOS8REjkAGC8/EjkvEjkvOS8SORE5LzkvMTABAyY1NDYzMhYXNjY3NjYzMhYVBwYHBgYHBgcOBBUUFhcWFQcGFRQXBgYVFxQjIiYnJiYnJicmJyYnJicGBwYHNCYnJicmJicmJyYnJjU3NycnNAE2Ab2HBi0YM5ZbKRODejgcJz0BCg0XFggECho5i0MZVkQrBQkFMxACCAcyFRMOEQ0HHx4NCQdmZ22MSQIVCQMDBgwJBQUODwIBAwQBAGYCdQIeGAwpO7fmHxGMhC5QIAgDAQMSGA4JGFTiWzAfS+tmPwcMEAgHDRoNFAsHHhoXCwUDCSUOBhINrlt6nEQVDx0ODgwGAwIOEQYHCAoICAsYASN1AAAAAAEAAAABAAAAAAAAXw889QA7CAAAAAAApWPHrgAAAACtlYR0///+ZQfUBmkAAAALAAAAAAAAAAAAAQAABmn+ZQAACCH//wAAB9QAAQAAAAAAAAAAAAAAAAAAAM0GAAEAAAAAAAYAAAACOQAAB8sAcgewAE0HywByB9cADQXAAC4GUACLBlIAPQZUACIFhQA4B64ASgeDAFUEZACEBtcAeAdKAIAHdwBIB0oAgAdKAEoHSgBoB0oAJAdKAEUHSgBgB0oAXwdK//8HSgAyB0oASAYUAEUGEgBHBggASAP0AEcEagATBEwATgSeAEkFiQA8BkoASwZOAEUGTgBFBlIASQZYAEwGWgBNBocATAaVAEwGUABABroAZQaVAEwGqgBWBocARQamAEgHYgBlBfQAPAXJACUF/gBIBlIARwZWAGAFjwBLBjUASAYlAEcGVgBIBhIARwWoAEAFqgBFBXUAGgWcACsGnABHBoUARwZQAEcGUABaBagAOQV/AEIFkQA8BYMAAgZKAD0GTABXBbQAVwZUAHsGSAA1BlQAMwb8AFMGFwAwBhgAMAYYADAGEgAvBhIALwcjADYHIwA2Bk4ATQZGAEkDgQA7ARsAOwI3ADsDUgA7AyMAcgMjAHIFWABNBVgATQMfAFMDHwA7AokALgKJAFMCNQAuAjUARgQSABUEEgAtA0gALwNIAEcB3wBHAd8ARwKsAGMCrABjBdsAswRaAHoEWgA5B0gASAVWAE0GFACcBhQAAQY1AEgEwgAYBY0APAUCAAIGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBycALQa0AEUIIQBNA6oAdAX8ANkHZABDBfwA+AdYADoHagBOB20AqAdtAKgGrABIBvwASQagABsHZABHB2QARwdWANMHcQBVB3MAVgO0AF0HEAAqBrAASQawAFMG8AB9BvAAfQWRAEsFkQBLBv4ATQb+AE0GFAAfB5EAMAYrAFcG6wA3BisAKQcbAL8HvAB0BxsAyQamAEcG/AA5B2oAqQfCAB4HWABTAAAAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgB1AHUAdQB1ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQE5ATkBOQABAAAAzQFSABAAAAAAAAIAEAATADgAAAH+//8ABgABAAAAFAD2AAEAAAAAAAAAEAAAAAEAAAAAAAEAFAAQAAEAAAAAAAIABwAkAAEAAAAAAAMACAArAAEAAAAAAAQAFAAzAAEAAAAAAAUADABHAAEAAAAAAAYAAABTAAEAAAAAAAcABwBTAAEAAAAAAAgABwBaAAEAAAAAAAkABwBhAAMAAQQJAAAAIABoAAMAAQQJAAEAKACIAAMAAQQJAAIADgCwAAMAAQQJAAMAEAC+AAMAAQQJAAQAKADOAAMAAQQJAAUAGAD2AAMAAQQJAAYAAAEOAAMAAQQJAAcADgEOAAMAAQQJAAgADgEcAAMAAQQJAAkADgEqT3JpZ2luYWwgbGljZW5jZUJFRk5PRytNb25vdHlwZVNvcnRzVW5rbm93bnVuaXF1ZUlEQkVGTk9HK01vbm90eXBlU29ydHNWZXJzaW9uIDAuMTFVbmtub3duVW5rbm93blVua25vd24ATwByAGkAZwBpAG4AYQBsACAAbABpAGMAZQBuAGMAZQBCAEUARgBOAE8ARwArAE0AbwBuAG8AdAB5AHAAZQBTAG8AcgB0AHMAVQBuAGsAbgBvAHcAbgB1AG4AaQBxAHUAZQBJAEQAQgBFAEYATgBPAEcAKwBNAG8AbgBvAHQAeQBwAGUAUwBvAHIAdABzAFYAZQByAHMAaQBvAG4AIAAwAC4AMQAxAFUAbgBrAG4AbwB3AG4AVQBuAGsAbgBvAHcAbgBVAG4AawBuAG8AdwBuAAAAAwAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAEEYACACmQAwApkAQAKZAFACmQAEACABpQAwAaUAQAGlAFABpQBwAaUABQCAAnMAsAJzQA0CAEZGAAAAEhEIQEgguAEDQE9IMiDeSDIg3EgyINpIMiDZSDIgrkgyIKFIMiCfSDIgj0gyIINIMiB+SDIgaEgyIGRIMiBgSDIgX0gyIF5IMiBdSDIgW0gyIFlIMiBVSDIguAHCskgyILgBwbJIMiC4AUCySDIguAE+skgyILgBPbJIMiC4AQSySDIguAECQJVIMiDdSDIg20gyILhIMiCiSDIgoEgyIJBIMiCOSDIghUgyIIRIMiCCSDIgfUgyIHhIMiB3SDIgaUgyIGVIMiBiSDIgWEgyEQkRCZCaB5CWB5CTB5CHB5B7B5B2B5ByB5BrB5BmB5BaB5BXB5BWByQIIgggCB4IHAgaCBgIFggUCBIIEAgOCAwICggICAYIBAgCCAAIAAFLsMBjAEtiILD2UyO4AQpRWrAFI0IBsBJLAEtUQrkAAQfAhY0WKysrKysrKysrKysrKysrKysrKxgrKysrKysrKysrKysBS1B5uQAfAdG2Bx/EBx9wBysrK0tTebkAkAHRtgeQxAeQcAcrKysYAbJQADJLYYtgHQArKysrKysrKysrKysrKysrKysrKysrKysBKysrKysrKysrKysrKysrKysrKysBRWlTQgFLUFixCABCWUNcWLEIAEJZswILChJDWGAbIVlCFhBwPrASQ1i5OyEYfhu6BAABqAALK1mwDCNCsA0jQrASQ1i5LUEtQRu6BAAEAAALK1mwDiNCsA8jQrASQ1i5GH47IRu6AagEAAALK1mwECNCsBEjQgFzc3MAAA==); }&#xA;@font-face { font-family: &quot;g_font_9&quot;; src: url(data:font/opentype;base64,AAEAAAANAIAAAwBQT1MvMmFqVnUAAADcAAAATmNtYXC/8yB+AAABLAAAADRjdnQgTw5I2QAAAWAAAAV0ZnBnbY+n6YkAAAbUAAAEI2dseWav/nuBAAAK+AAAAFRoZWFkuhmV8AAAC0wAAAA2aGhlYQ4+B1QAAAuEAAAAJGhtdHjKwDzQAAALqAAAAzRsb2NhELwQ5gAADtwAAAGcbWF4cAMrAWcAABB4AAAAIG5hbWW3qf4bAAAQmAAAAo5wb3N0AAMAAAAAEygAAAAgcHJlcG6IrVkAABNIAAACegAABAABkAAFAAAEAAQAAAAEAAQABAAAAAQAAGYCEgAAAQEBAQEBAQEBAQAAAAAAAAAAAAAAAAAAAAA/Pz8/AEAAIAAgCAACAADMBmkCmgAAAAAAAQADAAEAAAAMAAQAKAAAAAYABAABAAIAIOAA//8AAAAg4AD////jIAMAAQAAAAAAAAWRAAAFwQAABRsAWgWzAAQAAP/kAAAAAAEV/usAAAAABcEAAAAAAAD/5AAABaQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAD///////////////////////////////8AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA////////AAAAAAAyAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAADIAlQKZAEYARwEFAEAAdwBDACgAQQArAOYAOQCIAC8AJwC0AAMAKQAtAHoBRwAEAZQAYgXAAKwAxAKZArYAVQBaApkAKABCAIoAmQChAA0AKgBHAG4AcAW0ADYAPQBHAEcA/gGJAaQB6AJKAm4ABQAPACQAKgAqAIwAmACwANkA6wE5AT0BcgGRAZgBogHwBcAAHwA2ADsARwBHAFEAegC/AMIA5QI+AAgADgAWABYAJgBHAHEAswDZAOwBZwGIAcgB6QK2ADYAPABBAE4AUQBWAFoAiACVAJ0AsgC/AMMAxwDIANcBBwEpAUsBSwFxAYkBkgIWAlkCWQJaAnMCtwXwABYAGQAjACkAKgAqADEAPAA/AFEAUQBVAFsAdAB2AHkAgACXAKMAwQDKANwA8AEJAScBKwErATMBVAFrAWsBkQGrAcYB4QIkAioCQQJvAngCrgYXABEAJwArADEAPwBVAGEAYgBoAGkAbwBzAH8AfwCBAIQAhgCSAJcAmgCdAJ8AnwCrAK4AvQDPANIA3QDxAPIBDQElATMBOAFcAWgBfAGJAZwBnQGjAbYB0AHbAdsB/AIJAkMCkgOmBKgFFQWWBiIGtwbSABEAIAAyADwAPAA8AD0ARwBVAFYAVwBaAFsAXABcAHEAcwB0AHUAdgB8AIAAggCNAJ4AsQCyALIAsgC3AMQAxADRANkA3ADdAO8A8gD1APYBAQEDAQYBBwELARABFgEnAS4BMwE7AUoBTgFRAVUBWwFdAWQBaQFxAXIBkAGQAZQBmQGjAaYBpgGnAbEBswGzAbkBuwHGAccByAHaAfICGgIfAjUCNwI9AkkCUwJTAmMCdwKDAoYCkQKWApYClgLMAtAC0QLUAucC/AMJAygDNgM7A2QDdAOjA8sENwQ5BKAE1QTaBNwE3ATcBOkE/gUeBTgFWAWBBZYF2AXdBhMGZAaiBrYG1gbfBugG+geHAA0AJABDAFUAWgBuAHIAfQCKAIsAjwCXAKYAqQC2ALYAtwDEAM8A0wDaANsA5QDlAOsA7gELARUBHAEgAUYBRgFGAUkBWQFaAW0BcgF1AXYBfgGRAZIBnAGmAacBqQHBAcMBxQHeAd8B4QHyAfMB+QH9Af0CAAIVAhYCGQIaAh4CHwIiAi8CNAI0Aj0CSAJaAloCXQJkAm4CeAKBAoECiAKQAqYCqAKrAr8CwwLEAssC3ALgAvAC+wMLAw8DJgMrAzQDNQNcA3IDiwONA54DoAOkA60DxgPRA9ED2QP7BAAEUAR6BI4E2QUABQEFFQU2BV8FggWiBbkF5gXvBgsGFQYaBh0GMQZJBkoGVQZrBn4GlwbIBvYHAwcWBywHSQeHB8cAjwCdAI0AAAAAAAAAAAAAAAAAAAByAE0ApwBcAZsAKAArAAEAIgC5BFsAZQMeAoUBWQDCA/wAwgP8AJsBKAB+AL0BEgQ3AEsAqQErAH4BXwGYAEoAVwXAAJ0BZADHANoAfAA9ALIBvwAeAyYBOgDYAAIALQDZAJUBHAC/AgcCrgWOAakAiQA8APgARwA1AG4DvQPVA7sCWABrAPABrgEFADcB1ANcAW4BxwMKAmIC8ALaA1wBOAT+Be8FwQAAARgAPALtArIAtQAgApMCXgR9Ay5ANTQzMjEwLy4tLCsqKSgnJiUkIyIhIB8eHRwbGhkYFxYVFBMSERAPDg0MCwoJCAcGBQQDAgEALEUjRmAgsCZgsAQmI0hILSxFI0YjYSCwJmGwBCYjSEgtLEUjRmCwIGEgsEZgsAQmI0hILSxFI0YjYbAgYCCwJmGwIGGwBCYjSEgtLEUjRmCwQGEgsGZgsAQmI0hILSxFI0YjYbBAYCCwJmGwQGGwBCYjSEgtLAEQIDwAPC0sIEUjILDNRCMguAFaUVgjILCNRCNZILDtUVgjILBNRCNZILAEJlFYIyCwDUQjWSEhLSwgIEUYaEQgsAFgIEWwRnZoikVgRC0sAbELCkMjQ2UKLSwAsQoLQyNDCy0sALBGI3CxAUY+AbBGI3CxAkZFOrECAAgNLSxFsEojREWwSSNELSwgRbADJUVhZLBQUVhFRBshIVktLLABQ2MjYrAAI0KwDystLCBFsABDYEQtLAGwBkOwB0NlCi0sIGmwQGGwAIsgsSzAioy4EABiYCsMZCNkYVxYsANhWS0sRbARK7BHI0SwR3rkGC0suAGmVFiwCUO4AQBUWLkASv+AsUmARERZWS0sigNFioqHsBErsEcjRLBHeuQYLSwtLEtSWCFFRBsjRYwgsAMlRVJYRBshIVlZLSwBGC8tLCCwAyVFsEkjREWwSiNERWUjRSCwAyVgaiCwCSNCI2iKamBhILAairAAUnkhshpKQLn/4ABKRSCKVFgjIbA/GyNZYUQcsRQAilJ5s0lAIElFIIpUWCMhsD8bI1lhRC0ssRARQyNDCy0ssQ4PQyNDCy0ssQwNQyNDCy0ssQwNQyNDZQstLLEOD0MjQ2ULLSyxEBFDI0NlCy0sS1JYRUQbISFZLSwBILADJSNJsEBgsCBjILAAUlgjsAIlOCOwAiVlOACKYzgbISEhISFZAS0sRWmwCUNgihA6LSwBsAUlECMgivUAsAFgI+3sLSwBsAUlECMgivUAsAFhI+3sLSwBsAYlEPUA7ewtLCCwAWABECA8ADwtLCCwAWEBECA8ADwtLLArK7AqKi0sALAHQ7AGQwstLD6wKiotLDUtLHawSyNwECCwS0UgsABQWLABYVk6LxgtLCEhDGQjZIu4QABiLSwhsIBRWAxkI2SLuCAAYhuyAEAvK1mwAmAtLCGwwFFYDGQjZIu4FVViG7IAgC8rWbACYC0sDGQjZIu4QABiYCMhLSy0AAEAAAAVsAgmsAgmsAgmsAgmDxAWE0VoOrABFi0stAABAAAAFbAIJrAIJrAIJrAIJg8QFhNFaGU6sAEWLSxFIyBFILEEBSWKUFgmYYqLGyZgioxZRC0sRiNGYIqKRiMgRopgimG4/4BiIyAQI4qxS0uKcEVgILAAUFiwAWG4/8CLG7BAjFloATotLLAzK7AqKi0AAAIBAAAABQAFAAADAAcAKrUEkAAHkAG4AjSyAAoEvgE6AAAABQE6AAMCLwAAL/7lEOUAP/7lEOUxMCERIRElIREhAQAEAPwgA8D8QAUA+wAgBMAAAAEAAAABAAAAAAAAXw889QA7CAAAAAAApWPHrgAAAACtlYR0///+ZQfUBmkAAAALAAAAAAAAAAAAAQAABmn+ZQAACCH//wAAB9QAAQAAAAAAAAAAAAAAAAAAAM0GAAEAAAAAAAYAAAACOQAAB8sAcgewAE0HywByB9cADQXAAC4GUACLBlIAPQZUACIFhQA4B64ASgeDAFUEZACEBtcAeAdKAIAHdwBIB0oAgAdKAEoHSgBoB0oAJAdKAEUHSgBgB0oAXwdK//8HSgAyB0oASAYUAEUGEgBHBggASAP0AEcEagATBEwATgSeAEkFiQA8BkoASwZOAEUGTgBFBlIASQZYAEwGWgBNBocATAaVAEwGUABABroAZQaVAEwGqgBWBocARQamAEgHYgBlBfQAPAXJACUF/gBIBlIARwZWAGAFjwBLBjUASAYlAEcGVgBIBhIARwWoAEAFqgBFBXUAGgWcACsGnABHBoUARwZQAEcGUABaBagAOQV/AEIFkQA8BYMAAgZKAD0GTABXBbQAVwZUAHsGSAA1BlQAMwb8AFMGFwAwBhgAMAYYADAGEgAvBhIALwcjADYHIwA2Bk4ATQZGAEkDgQA7ARsAOwI3ADsDUgA7AyMAcgMjAHIFWABNBVgATQMfAFMDHwA7AokALgKJAFMCNQAuAjUARgQSABUEEgAtA0gALwNIAEcB3wBHAd8ARwKsAGMCrABjBdsAswRaAHoEWgA5B0gASAVWAE0GFACcBhQAAQY1AEgEwgAYBY0APAUCAAIGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBk4ARwZOAEcGTgBHBycALQa0AEUIIQBNA6oAdAX8ANkHZABDBfwA+AdYADoHagBOB20AqAdtAKgGrABIBvwASQagABsHZABHB2QARwdWANMHcQBVB3MAVgO0AF0HEAAqBrAASQawAFMG8AB9BvAAfQWRAEsFkQBLBv4ATQb+AE0GFAAfB5EAMAYrAFcG6wA3BisAKQcbAL8HvAB0BxsAyQamAEcG/AA5B2oAqQfCAB4HWABTAAAAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgAqACoAKgABAAAAzQFSABAAAAAAAAIAEAATADgAAAH+//8ABgABAAAAFAD2AAEAAAAAAAAAEAAAAAEAAAAAAAEAFAAQAAEAAAAAAAIABwAkAAEAAAAAAAMAFAArAAEAAAAAAAQAFAA/AAEAAAAAAAUADABTAAEAAAAAAAYAFABfAAEAAAAAAAcABwBzAAEAAAAAAAgABwB6AAEAAAAAAAkABwCBAAMAAQQJAAAAIACIAAMAAQQJAAEAKACoAAMAAQQJAAIADgDQAAMAAQQJAAMAKADeAAMAAQQJAAQAKAEGAAMAAQQJAAUAGAEuAAMAAQQJAAYAKAFGAAMAAQQJAAcADgFuAAMAAQQJAAgADgF8AAMAAQQJAAkADgGKT3JpZ2luYWwgbGljZW5jZUJFRk5PSCtNb25vdHlwZVNvcnRzVW5rbm93bkJFRk5PSCtNb25vdHlwZVNvcnRzQkVGTk9IK01vbm90eXBlU29ydHNWZXJzaW9uIDAuMTFCRUZOT0grTW9ub3R5cGVTb3J0c1Vua25vd25Vbmtub3duVW5rbm93bgBPAHIAaQBnAGkAbgBhAGwAIABsAGkAYwBlAG4AYwBlAEIARQBGAE4ATwBIACsATQBvAG4AbwB0AHkAcABlAFMAbwByAHQAcwBSAGUAZwB1AGwAYQByAEIARQBGAE4ATwBIACsATQBvAG4AbwB0AHkAcABlAFMAbwByAHQAcwBCAEUARgBOAE8ASAArAE0AbwBuAG8AdAB5AHAAZQBTAG8AcgB0AHMAVgBlAHIAcwBpAG8AbgAgADAALgAxADEAQgBFAEYATgBPAEgAKwBNAG8AbgBvAHQAeQBwAGUAUwBvAHIAdABzAFUAbgBrAG4AbwB3AG4AVQBuAGsAbgBvAHcAbgBVAG4AawBuAG8AdwBuAAAAAwAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAEEYACACmQAwApkAQAKZAFACmQAEACABpQAwAaUAQAGlAFABpQBwAaUABQCAAnMAsAJzQA0CAEZGAAAAEhEIQEgguAEDQE9IMiDeSDIg3EgyINpIMiDZSDIgrkgyIKFIMiCfSDIgj0gyIINIMiB+SDIgaEgyIGRIMiBgSDIgX0gyIF5IMiBdSDIgW0gyIFlIMiBVSDIguAHCskgyILgBwbJIMiC4AUCySDIguAE+skgyILgBPbJIMiC4AQSySDIguAECQJVIMiDdSDIg20gyILhIMiCiSDIgoEgyIJBIMiCOSDIghUgyIIRIMiCCSDIgfUgyIHhIMiB3SDIgaUgyIGVIMiBiSDIgWEgyEQkRCZCaB5CWB5CTB5CHB5B7B5B2B5ByB5BrB5BmB5BaB5BXB5BWByQIIgggCB4IHAgaCBgIFggUCBIIEAgOCAwICggICAYIBAgCCAAIAAFLsMBjAEtiILD2UyO4AQpRWrAFI0IBsBJLAEtUQrkAAQfAhY0WKysrKysrKysrKysrKysrKysrKxgrKysrKysrKysrKysBS1B5uQAfAdG2Bx/EBx9wBysrK0tTebkAkAHRtgeQxAeQcAcrKysYAbJQADJLYYtgHQArKysrKysrKysrKysrKysrKysrKysrKysBKysrKysrKysrKysrKysrKysrKysBRWlTQgFLUFixCABCWUNcWLEIAEJZswILChJDWGAbIVlCFhBwPrASQ1i5OyEYfhu6BAABqAALK1mwDCNCsA0jQrASQ1i5LUEtQRu6BAAEAAALK1mwDiNCsA8jQrASQ1i5GH47IRu6AagEAAALK1mwECNCsBEjQgFzc3MAAA==); }&#xA;</svg:style><svg:clipPath id="clippath3" transform="matrix(255.12 0 0 108.48 170.16 645.8604)"><svg:rect x="0" y="0" width="1063" height="452" clip-rule="nonzero"></svg:rect></svg:clipPath></svg:defs><svg:g transform=""><svg:text transform="matrix(10.9755 0 0 10.98 294.66 795.7403) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_3" font-size="1px" y="0"></svg:tspan><svg:tspan x="0" y="0" font-family="g_font_3" font-size="1px" fill="rgb(0,0,0)">3</svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="0" x="0.5576" fill="rgb(0,0,0)"> </svg:tspan></svg:text><svg:text transform="matrix(7.9767 0 0 7.98 49.62 38.6603) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_2" font-size="1px" y="0" x="0 0.7379 1.0164 1.7393 2.4622 3.0191 3.687 4.3549 4.6334 5.1903 5.7472 6.3112 6.8752 27.6433 28.2002 28.7571 29.314 29.8709 30.1498 30.7067 31.2636 31.5425 32.3764 32.6553 33.1562 33.4351 33.992 34.556" fill="rgb(0,0,0)">© UCLES 2019 0610/13/M/J/19 </svg:tspan></svg:text><svg:text transform="matrix(10.9755 0 0 10.98 491.28 38.6603) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_3" font-size="1px" y="0" x="0 0.3341 0.9462 1.5583 1.9484 2.5605 2.8395 3.4516 4.0087 4.5658" fill="rgb(0,0,0)">[Turn over</svg:tspan></svg:text><svg:text transform="matrix(7.9767 0 0 7.98 545.7 38.6603) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_2" font-size="1px" y="0" x="0" fill="rgb(0,0,0)"> </svg:tspan></svg:text><svg:text transform="matrix(10.9755 0 0 10.98 49.62 769.4603) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_3" font-size="1px" y="0" x="0 0.5575" fill="rgb(0,0,0)">3 </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="0" x="1.9407 2.5531 3.1105 3.6679 3.9469 4.5043 5.0617 5.6191 5.8985 6.4559 7.0133 7.3477 7.9051 8.4625 9.0199 9.2989 9.8003 10.3577 10.9151 11.6385 12.1399 12.4134 12.9708 13.5282 13.8072 14.3646 14.699 15.2564 15.8138 16.3712 16.5946 17.096 17.9304 18.2098" fill="rgb(0,0,0)">The photograph shows an organism. </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="1.153" x="0" fill="rgb(0,0,0)"> </svg:tspan></svg:text></svg:g><svg:g clip-path="url(#clippath3)"><svg:g transform="matrix(255.12 0 0 108.48 170.16 645.8604)"><svg:image xlink:href="data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAABCcAAAHECAIAAACFv9d4ABYA0UlEQVR4nAD//wAAAP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7u7u7////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////3d3d7u7u7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7u7u7u7u7t3d3czMzMzMzLu7u6qqqqqqqqqqqqqqqszMzN3d3f///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////u7u7u7u7u7u7u7u7u7u7d3d3d3d3MzMy7u7uqqqqqqqqIiIh3d3d3d3eIiIi7u7vd3d3u7u7////u7u7////u7u7u7u7////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u////7u7u7u7u7u7u7u7u3d3d3d3du7u7u7u7qqqqmZmZd3d3ZmZmd3d3iIiIu7u73d3d7u7u7u7u7u7u3d3d3d3d7u7u////////////////////////////////////////////////////////////7u7u////////////////////////////////////7u7u////////////////////////////////7u7u////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7v///////+7u7v///93d3d3d3czMzLu7u6qqqpmZmYiIiHd3d3d3d3d3d6qqqt3d3e7u7u7u7szMzLu7u7u7u8zMzN3d3e7u7u7u7u7u7v///////////////////////////////////////////////////////////+7u7u7u7v///////////+7u7u7u7u7u7v///+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7////u7u7////////////d3d3MzMzd3d3u7u7////u7u7////u7u7u7u7d3d3MzMzMzMy7u7uqqqqZmZmZmZmIiIiIiIiqqqrd3d3u7u7d3d27u7uqqqqZmZmZmZmZmZm7u7u7u7vMzMzd3d3u7u7u7u7////////u7u7////////////////u7u7////////////d3d3d3d3////////////u7u7u7u7u7u7////u7u7d3d3MzMzMzMzd3d3u7u7////////////////////////////////////////////u7u7////////////////u7u7u7u7MzMy7u7vMzMzd3d3d3d3d3d3u7u7u7u7////////////////////////u7u7////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u////////////////////////////////////7u7u7u7u7u7u////////3d3dqqqqmZmZ3d3d7u7u////7u7u7u7u////7u7u7u7u3d3d3d3dzMzMu7u7u7u7qqqqqqqqmZmZqqqq3d3d3d3d7u7uzMzMqqqqiIiId3d3d3d3iIiIiIiIiIiImZmZmZmZu7u77u7u7u7u////////////////7u7u7u7u7u7u////zMzMzMzM7u7u////////////7u7u7u7u3d3d7u7u3d3du7u7qqqqmZmZmZmZqqqqu7u73d3d////////7u7u////////////////////////////////////////////7u7uu7u7iIiId3d3d3d3mZmZqqqqmZmZqqqqu7u7zMzM3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////+7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzN3d3d3d3e7u7v///////////////////////+7u7u7u7u7u7t3d3e7u7u7u7t3d3aqqqru7u+7u7v///////////+7u7v///+7u7u7u7u7u7t3d3czMzMzMzMzMzLu7u7u7u6qqqqqqqru7u8zMzN3d3bu7u4iIiHd3d4iIiIiIiHd3d4iIiHd3d3d3d5mZmaqqqru7u8zMzO7u7v///////+7u7u7u7u7u7t3d3czMzMzMzO7u7u7u7v///////93d3d3d3e7u7u7u7u7u7t3d3bu7u5mZmWZmZmZmZmZmZoiIiLu7u93d3e7u7v///////+7u7v///////////+7u7u7u7u7u7u7u7v///////+7u7szMzJmZmXd3d3d3d4iIiHd3d3d3d3d3d4iIiIiIiKqqqru7u93d3f///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////u7u7d3d3d3d3d3d3MzMy7u7u7u7u7u7u7u7u7u7u7u7vMzMzd3d3u7u7////////////////////u7u7u7u7u7u7u7u7d3d3d3d2ZmZm7u7vd3d3u7u7////u7u7u7u7////u7u7////u7u7u7u7u7u7d3d3d3d3MzMzMzMy7u7uZmZmZmZmqqqq7u7u7u7uqqqqIiIiIiIh3d3eIiIiIiIiIiIiIiIiZmZmZmZmZmZmqqqrMzMzd3d3u7u7////////u7u7d3d3MzMzMzMzMzMzd3d3u7u7////u7u7d3d3d3d3u7u7u7u7u7u7u7u7MzMyqqqqIiIhmZmZmZmZ3d3eqqqq7u7vMzMzu7u7////////u7u7////u7u7d3d3MzMzMzMzu7u7////////////u7u7MzMyqqqqIiIiIiIh3d3dmZmZ3d3dmZmZ3d3d3d3eZmZm7u7vu7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u////////////////////7u7u////////////////////////////////7u7u////////////////////7u7u3d3d3d3dqqqqmZmZmZmZqqqqu7u7qqqqqqqqqqqqu7u7zMzM7u7u7u7u////////////////7u7u7u7u7u7u3d3du7u7iIiIiIiIu7u77u7u7u7u////////7u7u7u7u////7u7u////7u7u7u7u7u7u3d3d3d3dzMzMu7u7mZmZmZmZqqqqqqqqu7u7mZmZiIiIiIiIiIiIiIiImZmZmZmZmZmZqqqqqqqqmZmZqqqqqqqqzMzM3d3d////////7u7u7u7u3d3dzMzMu7u7u7u73d3d7u7u////7u7u////7u7u7u7u////7u7u3d3du7u7mZmZd3d3d3d3d3d3mZmZqqqqu7u7zMzM7u7u////7u7u////7u7u3d3dzMzMu7u73d3d7u7u////////////7u7u3d3du7u7qqqqmZmZiIiId3d3d3d3d3d3d3d3d3d3qqqqzMzM7u7u////////////////////////7u7u////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7t3d3d3d3czMzLu7u7u7u7u7u7u7u7u7u93d3d3d3e7u7v///////////+7u7u7u7t3d3e7u7u7u7v///////////////+7u7v///////////////////+7u7szMzLu7u6qqqqqqqqqqqqqqqqqqqru7u7u7u7u7u7u7u8zMzO7u7u7u7v///////////////+7u7u7u7t3d3bu7u4iIiIiIiJmZmd3d3f///+7u7u7u7v///+7u7u7u7u7u7v///////+7u7u7u7u7u7u7u7szMzLu7u7u7u5mZmYiIiIiIiKqqqoiIiHd3d4iIiJmZmZmZmaqqqqqqqqqqqqqqqpmZmaqqqpmZmZmZmaqqqru7u93d3e7u7v///+7u7u7u7t3d3aqqqqqqqru7u8zMzO7u7u7u7v///+7u7u7u7u7u7u7u7u7u7t3d3bu7u5mZmYiIiHd3d5mZmZmZmaqqqszMzN3d3e7u7u7u7u7u7u7u7u7u7ru7u6qqqru7u93d3f///////////////+7u7qqqqqqqqru7u6qqqpmZmXd3d3d3d3d3d2ZmZnd3d5mZmczMzO7u7u7u7v///+7u7v///////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3u7u7u7u7d3d3d3d3MzMy7u7uqqqqqqqqqqqqZmZmqqqqqqqrMzMzd3d3u7u7u7u7u7u7d3d3MzMy7u7vd3d3u7u7d3d3MzMzd3d3d3d3u7u7u7u7u7u7////u7u7u7u7u7u7d3d3d3d3d3d3MzMzMzMzMzMy7u7vMzMzMzMzMzMzMzMzd3d3d3d3u7u7////////////////u7u7u7u7d3d27u7uZmZmIiIiqqqrd3d3u7u7u7u7////u7u7////u7u7////u7u7u7u7u7u7u7u7u7u7d3d3d3d27u7uqqqqIiIiIiIiIiIiZmZmZmZmZmZmIiIiZmZmqqqqqqqq7u7uqqqqqqqqZmZmZmZmZmZmZmZmZmZmqqqrMzMzu7u7////////u7u7MzMzMzMyZmZmZmZmqqqq7u7vd3d3u7u7////u7u7u7u7u7u7u7u7d3d27u7uqqqqZmZmIiIiZmZmqqqq7u7vMzMzd3d3u7u7u7u7u7u7u7u7d3d2qqqqZmZmqqqrMzMzu7u7////////u7u67u7uZmZm7u7vMzMy7u7uqqqqZmZmIiIiIiIh3d3d3d3eZmZm7u7vd3d3u7u7////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u3d3d3d3dzMzM3d3dzMzMu7u7u7u7qqqqqqqqmZmZmZmZmZmZqqqqu7u73d3d3d3d3d3dzMzMqqqqmZmZu7u7u7u7zMzMzMzM3d3d7u7u7u7u7u7u7u7u////7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3dzMzM3d3dzMzM3d3dzMzM3d3d3d3d7u7u////////////7u7u7u7u3d3dzMzMmZmZiIiImZmZu7u77u7u////7u7u7u7u7u7u7u7u7u7u////7u7u7u7u3d3d3d3dzMzM3d3du7u7qqqqmZmZd3d3AP//AAB3d3eZmZmqqqqZmZmZmZmZmZmqqqq7u7u7u7u7u7u7u7uqqqqZmZmZmZmZmZmIiIiZmZm7u7vd3d3u7u7////u7u7u7u67u7uIiIh3d3d3d3eqqqrMzMzu7u7u7u7////u7u7u7u7u7u7d3d3MzMy7u7uqqqqZmZmZmZmZmZmqqqq7u7vMzMzd3d3u7u7////u7u7d3d27u7uIiIiIiIi7u7vd3d3///////////+7u7uZmZnMzMzd3d3d3d3MzMy7u7uZmZmZmZl3d3d3d3eIiIiZmZnMzMzu7u7////////u7u7u7u7u7u7////u7u7u7u7u7u7////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u3d3d7u7u3d3d3d3dzMzMzMzMu7u7u7u7u7u7qqqqqqqqmZmZqqqqqqqqzMzM3d3dzMzMzMzMmZmZmZmZqqqqzMzMu7u73d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u7u7u7u7u////7u7u7u7u7u7u3d3d3d3dzMzMzMzMzMzMzMzM3d3d3d3d3d3d7u7u////////7u7u7u7u3d3dzMzMqqqqd3d3d3d3mZmZ3d3d3d3d7u7u7u7u7u7u////7u7u7u7u7u7u3d3dzMzMzMzMzMzMzMzMzMzMu7u7iIiId3d3d3d3iIiImZmZqqqqmZmZmZmZqqqqu7u7zMzMzMzMu7u7zMzMqqqqqqqqmZmZmZmZmZmZu7u7u7u73d3d7u7u7u7u3d3dqqqqd3d3ZmZmZmZmiIiIqqqq3d3d////7u7u7u7u7u7u7u7u7u7u3d3d3d3du7u7u7u7mZmZmZmZmZmZmZmZu7u7zMzM3d3d////////3d3dmZmZZmZmZmZmiIiIzMzM7u7u////3d3dqqqqqqqq3d3d7u7u7u7u3d3dzMzMu7u7qqqqmZmZd3d3iIiImZmZzMzM3d3d////////7u7u7u7u3d3dzMzMzMzM3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////+7u7u7u7u7u7t3d3d3d3czMzMzMzMzMzLu7u7u7u7u7u6qqqqqqqqqqqru7u7u7u8zMzMzMzMzMzKqqqqqqqpmZmaqqqqqqqru7u93d3czMzO7u7u7u7v///+7u7v///+7u7u7u7v///+7u7v///+7u7u7u7u7u7u7u7t3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzO7u7u7u7v///+7u7u7u7t3d3czMzJmZmWZmZmZmZoiIiKqqqru7u93d3e7u7v///+7u7v///+7u7u7u7t3d3czMzLu7u7u7u8zMzMzMzLu7u4iIiIiIiIiIiJmZmaqqqqqqqqqqqqqqqqqqqqqqqru7u7u7u8zMzMzMzLu7u6qqqru7u6qqqqqqqpmZmbu7u8zMzN3d3d3d3czMzKqqqoiIiHd3d2ZmZnd3d5mZmczMzN3d3e7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3aqqqpmZmZmZmYiIiJmZmZmZmbu7u8zMzO7u7u7u7szMzJmZmXd3d2ZmZoiIiLu7u93d3f///93d3ZmZmbu7u93d3e7u7t3d3d3d3d3d3czMzKqqqpmZmYiIiHd3d4iIiLu7u93d3f///+7u7u7u7szMzLu7u6qqqpmZmd3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7////u7u7////u7u7u7u7d3d3d3d3d3d3MzMzMzMzMzMzMzMy7u7u7u7u7u7uqqqq7u7u7u7vMzMzd3d3MzMzMzMyqqqqqqqqZmZmIiIiZmZm7u7vMzMzu7u7////u7u7////////////u7u7////u7u7////u7u7u7u7u7u7u7u7d3d3MzMzMzMy7u7u7u7u7u7u7u7u7u7vMzMzd3d3u7u7u7u7u7u7d3d27u7uIiIhVVVVVVVVVVVVmZmaZmZnMzMzd3d3////u7u7u7u7u7u7d3d3d3d3MzMy7u7u7u7vMzMy7u7uqqqqZmZmIiIiZmZmqqqqqqqqZmZmZmZmqqqqqqqq7u7u7u7u7u7vMzMzMzMy7u7vMzMzMzMyqqqqqqqqZmZmZmZmqqqrMzMzd3d27u7uqqqqZmZmIiIh3d3dmZmaIiIiqqqrMzMzd3d3d3d3d3d3u7u7u7u7d3d3d3d3MzMzMzMyqqqqZmZmIiIiIiIiIiIiZmZmqqqrd3d3d3d3d3d27u7uZmZmIiIiIiIiZmZnMzMzd3d27u7uZmZnMzMzd3d3d3d3d3d3MzMzMzMy7u7uqqqqZmZmIiIh3d3d3d3eqqqrd3d3////u7u7d3d3MzMy7u7uqqqqqqqq7u7vd3d3u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////7u7u7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3dzMzMu7u7u7u7u7u7u7u7zMzM3d3d3d3d3d3dzMzMu7u7mZmZZmZmd3d3mZmZ3d3d7u7u////////7u7u////////7u7u////7u7u////7u7u7u7u7u7u7u7u3d3d3d3dzMzMu7u7u7u7qqqqqqqqqqqqu7u7zMzM3d3d7u7u7u7u3d3dzMzMiIiIZmZmVVVVVVVVVVVVZmZmmZmZzMzM7u7u7u7u7u7u7u7u3d3d3d3dzMzMu7u7zMzMzMzMu7u7u7u7u7u7mZmZmZmZmZmZqqqqqqqqmZmZqqqqqqqqqqqqqqqqu7u7u7u7zMzMzMzMzMzMu7u7u7u7qqqqmZmZiIiImZmZu7u73d3dzMzMu7u7mZmZmZmZiIiId3d3d3d3iIiIqqqqmZmZiIiIqqqq7u7u3d3d7u7u7u7u3d3d3d3du7u7qqqqmZmZiIiIiIiIiIiImZmZzMzM3d3d3d3dzMzMqqqqmZmZiIiIiIiIqqqqu7u7mZmZmZmZu7u73d3dzMzMzMzM3d3dzMzMu7u7u7u7qqqqiIiId3d3d3d3qqqqzMzM3d3d7u7uzMzMu7u7qqqqmZmZiIiIiIiImZmZzMzM3d3d7u7u////7u7u////////7u7u////////////////////////////////////7u7u////////////7u7u////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////+7u7v///////////////////////////////+7u7u7u7u7u7u7u7u7u7u7u7v///+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3bu7u7u7u6qqqru7u8zMzN3d3d3d3d3d3czMzJmZmXd3d2ZmZoiIiLu7u93d3f///////+7u7v///+7u7v///+7u7v///+7u7u7u7u7u7u7u7u7u7t3d3d3d3czMzLu7u7u7u7u7u5mZmZmZmZmZmaqqqt3d3d3d3e7u7t3d3czMzJmZmZmZmXd3d2ZmZlVVVWZmZoiIiKqqqszMzN3d3d3d3e7u7u7u7t3d3czMzMzMzN3d3d3d3czMzLu7u6qqqqqqqpmZmZmZmZmZmZmZmZmZmaqqqqqqqqqqqru7u7u7u7u7u7u7u8zMzMzMzMzMzLu7u6qqqpmZmYiIiIiIiKqqqszMzMzMzLu7u6qqqpmZmZmZmZmZmYiIiHd3d2ZmZkRERGZmZru7u93d3e7u7u7u7t3d3d3d3czMzMzMzLu7u7u7u5mZmYiIiIiIiJmZmbu7u93d3e7u7szMzLu7u6qqqoiIiIiIiIiIiHd3d2ZmZpmZmZmZmZmZmZmZmczMzMzMzMzMzMzMzMzMzKqqqpmZmYiIiIiIiJmZmbu7u8zMzMzMzLu7u6qqqpmZmYiIiHd3d2ZmZnd3d5mZmaqqqszMzN3d3e7u7v///////////////////////////+7u7v///////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////u7u7////////////////////////////u7u7////////////////u7u7////u7u7////u7u7////////////////////////u7u7u7u7////u7u7u7u7////u7u7////////////u7u7////u7u7u7u7u7u7u7u7d3d3MzMy7u7uqqqqqqqqqqqrMzMzd3d3u7u7u7u7MzMy7u7uZmZl3d3eIiIiqqqrd3d3u7u7u7u7////u7u7u7u7////u7u7////u7u7u7u7u7u7u7u7d3d3d3d3MzMzMzMzMzMy7u7u7u7uZmZmIiIiZmZmqqqq7u7vd3d3d3d3MzMy7u7uqqqqqqqqZmZmIiIh3d3dmZmZmZmaIiIiZmZnMzMzd3d3d3d3d3d3d3d3d3d3MzMy7u7vMzMy7u7uqqqqqqqqIiIiIiIiIiIiIiIiIiIiZmZmZmZmZmZmqqqqqqqq7u7u7u7vMzMzMzMzd3d3MzMy7u7uqqqqIiIh3d3eIiIiZmZm7u7u7u7uqqqqqqqqZmZmqqqqqqqqZmZmIiIh3d3dmZmZ3d3e7u7vd3d3u7u7d3d3d3d3MzMzMzMzMzMy7u7u7u7uqqqqZmZmZmZmZmZmqqqrMzMzd3d3d3d27u7uqqqqZmZmZmZmIiIh3d3dmZmZ3d3dmZmZmZmaZmZm7u7vMzMzd3d3d3d27u7uqqqqZmZmIiIiZmZmZmZmqqqrMzMy7u7uqqqqZmZmIiIh3d3d3d3dmZmZmZmZmZmZ3d3eIiIiqqqrMzMzu7u7////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////7u7u////7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3d7u7u////////////////////////7u7u7u7uzMzMzMzMzMzM7u7u7u7u////////////////////////7u7u////7u7u////7u7u////////7u7u////7u7u7u7u7u7u3d3d3d3d3d3d3d3dzMzMqqqqmZmZiIiIqqqqu7u7zMzM7u7u7u7u3d3dzMzMmZmZd3d3ZmZmmZmZzMzM7u7u7u7u////////7u7u////7u7u7u7u7u7u7u7u3d3d3d3d3d3dzMzMzMzMzMzM3d3du7u7u7u7qqqqmZmZd3d3mZmZu7u7zMzMzMzMzMzMu7u7qqqqu7u7qqqqiIiId3d3ZmZmZmZmd3d3mZmZqqqqu7u7zMzMzMzM3d3dzMzMzMzMu7u7zMzMqqqqiIiIZmZmZmZmZmZmZmZmd3d3d3d3iIiIiIiImZmZmZmZmZmZu7u7u7u7u7u7u7u7zMzMu7u7qqqqiIiId3d3ZmZmZmZmiIiIqqqqu7u7zMzMqqqqmZmZqqqqmZmZqqqqmZmZd3d3ZmZmd3d3qqqq3d3d3d3dzMzMzMzMu7u7zMzMu7u7u7u7u7u7qqqqmZmZiIiIiIiImZmZu7u7zMzMzMzMu7u7qqqqmZmZmZmZd3d3d3d3ZmZmVVVVZmZmZmZmiIiIqqqqzMzMzMzMzMzMzMzMu7u7qqqqqqqqmZmZmZmZqqqqqqqqqqqqqqqqmZmZmZmZd3d3d3d3ZmZmVVVVVVVVVVVVd3d3mZmZqqqqzMzM3d3d////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7t3d3czMzMzMzKqqqqqqqqqqqru7u93d3e7u7u7u7v///////////93d3czMzKqqqqqqqqqqqszMzN3d3e7u7v///////////////////////////////////////////////+7u7v///+7u7u7u7t3d3czMzLu7u7u7u7u7u6qqqqqqqpmZmZmZmYiIiJmZmczMzN3d3d3d3d3d3czMzKqqqoiIiGZmZnd3d5mZmczMzN3d3e7u7u7u7u7u7v///+7u7u7u7t3d3e7u7t3d3czMzMzMzMzMzMzMzMzMzMzMzN3d3bu7u7u7u5mZmYiIiIiIiKqqqru7u7u7u7u7u7u7u5mZmaqqqpmZmYiIiHd3d3d3d3d3d4iIiJmZmZmZmaqqqqqqqszMzLu7u8zMzMzMzMzMzLu7u6qqqoiIiGZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZoiIiJmZmaqqqru7u7u7u7u7u6qqqqqqqqqqqoiIiIiIiHd3d2ZmZmZmZnd3d5mZmczMzMzMzKqqqqqqqpmZmZmZmaqqqpmZmYiIiHd3d3d3d5mZmbu7u8zMzMzMzMzMzMzMzMzMzMzMzN3d3bu7u7u7u5mZmZmZmYiIiJmZmaqqqszMzMzMzN3d3czMzLu7u5mZmZmZmZmZmXd3d4iIiIiIiIiIiIiIiKqqqszMzN3d3d3d3d3d3czMzMzMzKqqqqqqqpmZmaqqqqqqqru7u8zMzLu7u6qqqoiIiIiIiHd3d2ZmZmZmZmZmZmZmZnd3d5mZmaqqqru7u93d3e7u7v///////////+7u7v///////////+7u7v///////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////u7u7u7u7u7u7d3d3MzMy7u7uZmZmZmZmqqqqqqqrMzMzd3d3u7u7u7u7////////u7u7d3d3MzMyqqqqqqqq7u7vMzMzd3d3u7u7////////////u7u7////////////////u7u7////u7u7u7u7d3d3d3d3d3d3MzMy7u7uqqqqZmZmZmZmqqqqqqqqZmZmZmZmIiIiZmZm7u7vd3d3d3d3d3d3MzMyqqqp3d3dVVVVVVVV3d3eqqqq7u7vd3d3u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3MzMy7u7uqqqrMzMzMzMzMzMzMzMy7u7vMzMyZmZmIiIiIiIiqqqq7u7vMzMzMzMyqqqqqqqqqqqqqqqqIiIiIiIh3d3eZmZmqqqq7u7uqqqq7u7u7u7u7u7vMzMy7u7vMzMzMzMzMzMy7u7uqqqp3d3d3d3dmZmZERERVVVVVVVVmZmZ3d3eIiIiqqqqqqqqqqqq7u7uqqqqqqqqqqqqZmZmZmZmIiIiIiIhmZmZmZmZ3d3eZmZnd3d3MzMzMzMyqqqqZmZmIiIiZmZmZmZmqqqqZmZmIiIiIiIiqqqrd3d3MzMzd3d3d3d3d3d3MzMzMzMzMzMy7u7u7u7uqqqqZmZmZmZmqqqrMzMzd3d3d3d27u7uqqqqqqqqqqqqqqqqIiIiZmZmZmZmZmZmZmZmqqqrMzMzd3d3d3d3d3d3MzMy7u7u7u7uqqqqqqqqZmZm7u7vMzMzMzMyqqqqqqqqIiIiIiIh3d3dmZmZmZmZmZmZmZmZmZmZ3d3eZmZmqqqq7u7vd3d3u7u7////u7u7////u7u7////////////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u////////////////////7u7u7u7u3d3d3d3dzMzMzMzMu7u7u7u7u7u7u7u7zMzM3d3d3d3d7u7u////////////7u7uzMzMqqqqu7u7u7u7zMzMzMzM3d3d7u7u////////////7u7u////////////7u7u7u7u3d3d3d3dzMzMzMzMzMzMu7u7u7u7u7u7qqqqmZmZmZmZiIiImZmZmZmZiIiImZmZqqqq3d3d3d3d3d3d3d3du7u7iIiIZmZmZmZmZmZmiIiIqqqqzMzM3d3d3d3d7u7u7u7u7u7u7u7u3d3dzMzMu7u7u7u7u7u7u7u7zMzMzMzMzMzM3d3dzMzMu7u7qqqqmZmZqqqqqqqqzMzMzMzMu7u7qqqqmZmZqqqqmZmZiIiIiIiImZmZmZmZu7u7zMzMzMzMzMzMu7u7zMzMzMzMu7u7u7u7zMzMzMzMu7u7qqqqmZmZd3d3VVVVVVVVZmZmiIiId3d3iIiIqqqqqqqqu7u7u7u7u7u7mZmZqqqqmZmZmZmZmZmZiIiId3d3ZmZmd3d3qqqqu7u73d3d3d3du7u7mZmZiIiIiIiIiIiImZmZmZmZmZmZiIiIqqqqzMzM3d3d3d3d3d3d3d3d3d3dzMzMzMzMu7u7u7u7qqqqmZmZmZmZqqqqzMzM3d3dzMzMu7u7qqqqqqqqqqqqqqqqmZmZiIiImZmZmZmZmZmZu7u7zMzM3d3d3d3d3d3dzMzMqqqqmZmZmZmZmZmZmZmZqqqqzMzMzMzMu7u7qqqqmZmZmZmZmZmZiIiIZmZmZmZmZmZmVVVVZmZmd3d3mZmZu7u7zMzM7u7u7u7u////////7u7u////////7u7u////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7v///+7u7v///////+7u7u7u7u7u7u7u7u7u7t3d3d3d3czMzLu7u7u7u7u7u7u7u7u7u8zMzN3d3d3d3e7u7v///////+7u7t3d3czMzMzMzMzMzMzMzMzMzN3d3e7u7v///////////+7u7v///////93d3d3d3bu7u7u7u7u7u8zMzLu7u7u7u8zMzLu7u7u7u7u7u7u7u5mZmYiIiJmZmYiIiIiIiIiIiJmZmd3d3d3d3d3d3e7u7szMzLu7u4iIiIiIiIiIiIiIiKqqqqqqqszMzMzMzN3d3e7u7u7u7u7u7t3d3czMzMzMzLu7u7u7u7u7u7u7u8zMzMzMzMzMzMzMzKqqqqqqqoiIiJmZmaqqqszMzMzMzMzMzKqqqpmZmZmZmYiIiIiIiIiIiIiIiJmZmczMzN3d3d3d3d3d3d3d3d3d3czMzLu7u7u7u7u7u8zMzLu7u7u7u6qqqnd3d3d3d3d3d4iIiHd3d5mZmaqqqqqqqpmZmZmZmaqqqqqqqqqqqpmZmZmZmYiIiJmZmZmZmYiIiGZmZmZmZoiIiKqqqt3d3czMzMzMzKqqqoiIiIiIiIiIiJmZmZmZmZmZmZmZmaqqqru7u8zMzN3d3d3d3d3d3d3d3d3d3czMzMzMzLu7u5mZmZmZmYiIiJmZmbu7u8zMzN3d3czMzLu7u6qqqqqqqqqqqoiIiIiIiJmZmaqqqqqqqqqqqru7u93d3d3d3d3d3czMzKqqqpmZmYiIiIiIiIiIiKqqqszMzMzMzN3d3czMzKqqqqqqqpmZmZmZmYiIiHd3d1VVVVVVVVVVVXd3d4iIiJmZmaqqqt3d3e7u7u7u7u7u7t3d3d3d3e7u7u7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////u7u7////////////u7u7////////////////////////////////////////u7u7////////u7u7////////////////////////u7u7u7u7u7u7////u7u7////u7u7////u7u7u7u7u7u7d3d27u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7vMzMzd3d3d3d3u7u7////u7u7u7u7d3d3d3d3d3d3d3d3MzMy7u7u7u7vu7u7u7u7////////d3d27u7uZmZl3d3d3d3eIiIiZmZm7u7vMzMy7u7u7u7u7u7uqqqq7u7u7u7uqqqqqqqqZmZmIiIh3d3d3d3eZmZm7u7vd3d3u7u7u7u7d3d3MzMyqqqqqqqqZmZmqqqq7u7vMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMy7u7vMzMy7u7u7u7u7u7uqqqqqqqqqqqqqqqqZmZmIiIh3d3eIiIiqqqrMzMy7u7uZmZmIiIiIiIh3d3eIiIiIiIiZmZmqqqq7u7vd3d3u7u7u7u7d3d3d3d3MzMy7u7uqqqqqqqq7u7vMzMzMzMyqqqqIiIiIiIh3d3eIiIiIiIiZmZmZmZmZmZmIiIiIiIiZmZmZmZmqqqqZmZmZmZmZmZmZmZmZmZl3d3d3d3dmZmZ3d3eIiIi7u7vd3d3d3d2qqqqZmZmZmZmIiIiIiIiZmZmZmZmIiIiIiIiZmZm7u7vd3d3d3d3u7u7d3d3d3d3d3d3d3d27u7uqqqqIiIiIiIiIiIiqqqrMzMzd3d3MzMy7u7uqqqqqqqqIiIh3d3eZmZmZmZm7u7u7u7u7u7u7u7vMzMzd3d3d3d3MzMy7u7uqqqqZmZmIiIh3d3eqqqrMzMzMzMzu7u7d3d3MzMy7u7uqqqqZmZmIiIh3d3dVVVVmZmZmZmZmZmZ3d3eIiIiZmZmqqqrd3d3u7u7d3d3d3d3d3d3MzMzd3d3d3d3////////////////////////////////u7u7////////u7u7////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////7u7u////7u7u////7u7u7u7u7u7u7u7u3d3du7u7qqqqqqqqmZmZqqqqqqqqqqqqqqqqu7u7u7u7zMzMzMzM3d3d3d3d7u7u////7u7u3d3d3d3d3d3dzMzMu7u7qqqqqqqq3d3d7u7uzMzMu7u7iIiId3d3ZmZmVVVVVVVVZmZmiIiIu7u7u7u7u7u7u7u7qqqqqqqqu7u7u7u7u7u7u7u7qqqqmZmZiIiId3d3iIiIqqqq3d3d7u7u3d3d3d3dzMzMu7u7u7u7qqqqu7u7zMzM3d3d3d3d7u7u3d3d3d3d7u7u3d3d3d3d3d3d3d3dzMzMu7u7u7u7u7u7qqqqmZmZqqqqqqqqmZmZmZmZd3d3d3d3d3d3qqqqu7u7qqqqmZmZd3d3d3d3d3d3iIiImZmZmZmZqqqqu7u73d3d7u7u3d3d7u7u3d3d3d3du7u7u7u7zMzMzMzMu7u7u7u7u7u7mZmZd3d3iIiImZmZiIiImZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZqqqqqqqqmZmZiIiIiIiIiIiId3d3ZmZmZmZmd3d3qqqq3d3d3d3du7u7qqqqmZmZiIiIiIiImZmZmZmZmZmZiIiIiIiIu7u7zMzM3d3d7u7u3d3d3d3d3d3dzMzMu7u7iIiId3d3d3d3d3d3qqqqu7u73d3d3d3dzMzMqqqqiIiIiIiIiIiIiIiIqqqqu7u7u7u7u7u7zMzMzMzMzMzMzMzMzMzMu7u7qqqqmZmZiIiIiIiImZmZu7u7zMzM3d3d3d3dzMzMu7u7qqqqqqqqiIiId3d3d3d3ZmZmd3d3d3d3d3d3d3d3mZmZqqqqu7u73d3d3d3d3d3d3d3dzMzM3d3dzMzM7u7u7u7u7u7u////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7v///////////+7u7u7u7v///+7u7t3d3bu7u7u7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqru7u7u7u7u7u7u7u8zMzN3d3d3d3e7u7u7u7u7u7u7u7t3d3czMzKqqqpmZmZmZmaqqqpmZmZmZmYiIiHd3d1VVVVVVVVVVVURERGZmZnd3d5mZmaqqqszMzLu7u8zMzMzMzLu7u7u7u7u7u8zMzLu7u6qqqoiIiHd3d4iIiKqqqt3d3d3d3e7u7szMzMzMzKqqqru7u7u7u7u7u8zMzN3d3d3d3e7u7u7u7u7u7u7u7u7u7t3d3d3d3czMzMzMzMzMzMzMzLu7u6qqqqqqqqqqqqqqqqqqqpmZmXd3d2ZmZmZmZoiIiLu7u8zMzKqqqnd3d3d3d3d3d3d3d4iIiIiIiJmZmbu7u8zMzN3d3e7u7t3d3d3d3czMzLu7u6qqqqqqqru7u7u7u7u7u6qqqpmZmYiIiIiIiIiIiIiIiJmZmaqqqqqqqpmZmaqqqpmZmZmZmYiIiKqqqqqqqpmZmZmZmZmZmZmZmYiIiGZmZmZmZnd3d6qqqszMzN3d3czMzLu7u5mZmZmZmYiIiJmZmZmZmaqqqpmZmYiIiJmZmbu7u93d3d3d3d3d3d3d3czMzMzMzKqqqpmZmXd3d2ZmZnd3d5mZmczMzO7u7t3d3czMzKqqqoiIiIiIiHd3d3d3d4iIiKqqqru7u7u7u7u7u6qqqru7u7u7u8zMzN3d3bu7u6qqqpmZmYiIiIiIiJmZmczMzN3d3czMzN3d3bu7u6qqqqqqqpmZmYiIiHd3d1VVVWZmZoiIiHd3d3d3d2ZmZoiIiKqqqru7u93d3d3d3e7u7t3d3d3d3czMzLu7u7u7u93d3f///+7u7t3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////u7u7////u7u7////u7u7u7u7u7u7u7u7u7u7u7u67u7u7u7uqqqqZmZmqqqqqqqqZmZmqqqqZmZmqqqqqqqq7u7u7u7u7u7u7u7vMzMzd3d3d3d3d3d3d3d3d3d3d3d3MzMy7u7uZmZmqqqqIiIiIiIiZmZmIiIhmZmZVVVVVVVVVVVVmZmZ3d3dmZmaqqqq7u7vMzMy7u7vMzMzMzMy7u7u7u7vMzMzMzMy7u7uqqqqZmZmIiIh3d3eZmZnMzMzd3d3d3d3d3d3MzMy7u7uqqqq7u7uqqqq7u7u7u7vMzMzd3d3d3d3u7u7d3d3d3d3MzMzMzMzMzMy7u7vMzMzMzMy7u7u7u7u7u7u7u7u7u7uqqqqqqqp3d3dmZmZmZmaIiIiqqqrMzMy7u7uIiIiIiIh3d3d3d3d3d3d3d3eIiIiZmZm7u7vMzMzd3d3d3d3d3d27u7uqqqqqqqqqqqq7u7vMzMy7u7u7u7uZmZmIiIiIiIiIiIiIiIiZmZmZmZmqqqq7u7uZmZmIiIiIiIiIiIiZmZmqqqqZmZmZmZmqqqqqqqqZmZl3d3dmZmZ3d3eqqqq7u7vMzMzd3d27u7uZmZmIiIiIiIiIiIiZmZm7u7uqqqqIiIiZmZmZmZm7u7vMzMzd3d27u7u7u7u7u7uqqqqZmZmIiIh3d3d3d3eZmZm7u7vd3d3d3d3MzMyqqqqIiIh3d3dmZmZmZmZmZmZ3d3eIiIiIiIiZmZmIiIiIiIiqqqq7u7vd3d3MzMy7u7uZmZl3d3d3d3eZmZmqqqrMzMzd3d3d3d27u7uqqqqZmZmZmZmZmZl3d3dmZmZ3d3eIiIiIiIh3d3dmZmZ3d3eZmZm7u7vMzMzu7u7u7u7u7u7d3d3MzMyqqqqZmZnMzMzd3d3d3d27u7vMzMzd3d3u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3d7u7u3d3d7u7u7u7u7u7u////////////////////////////////////////7u7u////7u7u7u7u////////////////////////////////////////////////7u7u////////7u7u////7u7u7u7u7u7uzMzMqqqqqqqqqqqqqqqqqqqqmZmZmZmZmZmZmZmZmZmZqqqqqqqqu7u7zMzMu7u7u7u7zMzMzMzM3d3d3d3d3d3d3d3dzMzMqqqqqqqqmZmZiIiImZmZqqqqqqqqiIiIZmZmVVVVZmZmZmZmZmZmiIiIu7u7u7u7u7u7u7u7u7u7zMzMu7u7u7u7u7u7qqqqu7u7u7u7qqqqiIiIiIiImZmZu7u73d3d3d3dzMzMzMzMu7u7u7u7qqqqmZmZqqqqu7u7u7u7zMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7zMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7qqqqmZmZiIiIZmZmVVVViIiIqqqqu7u7qqqqiIiIiIiId3d3ZmZmZmZmd3d3d3d3mZmZqqqqu7u7u7u7zMzMzMzMzMzMqqqqu7u7zMzMzMzMzMzMu7u7u7u7qqqqmZmZiIiIiIiIiIiImZmZqqqqmZmZiIiIiIiId3d3iIiIiIiIiIiImZmZmZmZqqqqmZmZmZmZqqqqiIiIZmZmd3d3mZmZqqqqu7u7zMzMu7u7qqqqiIiId3d3d3d3mZmZu7u7u7u7mZmZiIiIiIiImZmZu7u7u7u7u7u7qqqqqqqqqqqqmZmZiIiId3d3d3d3iIiIu7u7zMzM3d3du7u7qqqqiIiId3d3ZmZmVVVVVVVVZmZmZmZmiIiIiIiId3d3ZmZmiIiIqqqqzMzMu7u7u7u7qqqqiIiId3d3iIiIqqqqu7u73d3d3d3du7u7qqqqmZmZmZmZmZmZiIiIZmZmZmZmiIiImZmZiIiIiIiId3d3iIiIqqqqzMzM3d3d7u7u7u7u3d3du7u7iIiIiIiImZmZqqqqu7u7qqqqmZmZu7u7zMzM7u7u////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////93d3czMzN3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3e7u7u7u7u7u7v///////////+7u7u7u7u7u7t3d3e7u7t3d3f///////////////////////////////+7u7v///+7u7u7u7v///+7u7v///////+7u7t3d3bu7u7u7u7u7u6qqqqqqqqqqqpmZmZmZmYiIiJmZmZmZmZmZmZmZmbu7u7u7u7u7u7u7u7u7u7u7u7u7u8zMzN3d3d3d3czMzLu7u6qqqqqqqpmZmYiIiKqqqqqqqru7u6qqqoiIiGZmZmZmZlVVVWZmZoiIiKqqqqqqqru7u6qqqru7u8zMzLu7u7u7u7u7u7u7u7u7u7u7u6qqqpmZmZmZmZmZmbu7u8zMzMzMzN3d3czMzMzMzKqqqpmZmZmZmaqqqqqqqru7u7u7u7u7u7u7u7u7u8zMzMzMzLu7u8zMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u6qqqqqqqpmZmXd3d2ZmZmZmZnd3d6qqqru7u6qqqoiIiGZmZmZmZlVVVWZmZnd3d2ZmZoiIiKqqqqqqqqqqqru7u8zMzKqqqqqqqru7u8zMzMzMzLu7u7u7u7u7u6qqqpmZmYiIiIiIiJmZmaqqqqqqqoiIiHd3d3d3d2ZmZnd3d2ZmZoiIiIiIiJmZmZmZmZmZmaqqqqqqqoiIiHd3d2ZmZoiIiJmZmbu7u8zMzLu7u6qqqoiIiIiIiIiIiIiIiKqqqru7u5mZmXd3d2ZmZnd3d5mZmbu7u6qqqqqqqqqqqqqqqpmZmZmZmZmZmXd3d4iIiKqqqszMzN3d3bu7u5mZmXd3d2ZmZmZmZlVVVVVVVVVVVVVVVWZmZlVVVVVVVWZmZnd3d4iIiKqqqru7u7u7u6qqqoiIiHd3d4iIiKqqqru7u8zMzMzMzLu7u6qqqpmZmZmZmZmZmYiIiHd3d2ZmZnd3d5mZmZmZmZmZmYiIiHd3d5mZmbu7u+7u7u7u7u7u7ru7u4iIiHd3d2ZmZnd3d5mZmZmZmZmZmZmZmZmZmbu7u+7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u67u7u7u7vMzMzMzMzMzMzMzMy7u7u7u7uqqqqZmZmZmZmZmZmqqqrMzMzMzMzd3d3u7u7////u7u7u7u7d3d3MzMy7u7u7u7vu7u7u7u7u7u7////////////////////////////u7u7u7u7u7u7////u7u7u7u7d3d3MzMyqqqq7u7u7u7uqqqqqqqqqqqqqqqqqqqqqqqqZmZmIiIiZmZmZmZmZmZmqqqqqqqq7u7u7u7uqqqqqqqq7u7vMzMzd3d3MzMy7u7uqqqqZmZmZmZmIiIiIiIiZmZm7u7vMzMy7u7uqqqqIiIhmZmZmZmZ3d3eZmZmqqqqqqqq7u7u7u7vMzMzMzMzMzMy7u7u7u7u7u7u7u7uqqqqqqqqIiIiIiIiZmZmqqqrMzMzMzMzMzMzMzMyqqqqqqqqZmZmqqqqZmZmqqqqqqqqqqqqZmZmqqqqqqqq7u7u7u7vMzMzMzMzMzMzMzMzd3d3MzMy7u7u7u7u7u7u7u7uZmZl3d3dmZmZmZmZmZmaZmZm7u7u7u7uZmZl3d3d3d3dVVVVmZmZmZmZmZmZ3d3eIiIiZmZmZmZm7u7vMzMy7u7uqqqq7u7u7u7u7u7uqqqqqqqq7u7uZmZmZmZmIiIh3d3eIiIiqqqq7u7uqqqqIiIhmZmZmZmZmZmZ3d3d3d3eIiIiZmZmZmZmZmZm7u7uqqqqZmZlmZmZmZmZ3d3eZmZm7u7vMzMzMzMy7u7uqqqqZmZmIiIiZmZmqqqq7u7uZmZmIiIhmZmZ3d3eIiIi7u7u7u7vMzMy7u7u7u7u7u7uqqqqZmZl3d3d3d3eZmZmqqqrMzMy7u7uqqqqIiIh3d3d3d3dmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZ3d3eZmZmqqqqZmZmIiIh3d3eIiIiZmZmqqqrMzMzMzMy7u7uqqqqZmZmZmZmZmZmZmZl3d3d3d3eIiIiqqqq7u7uqqqqIiIh3d3eIiIi7u7vd3d3u7u7d3d27u7t3d3dmZmZmZmZ3d3eIiIiIiIiZmZmIiIiIiIiqqqrMzMzu7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////3d3du7u7u7u7u7u7zMzMzMzMu7u7u7u7qqqqmZmZiIiIiIiId3d3d3d3iIiIiIiIqqqqzMzM3d3d3d3d3d3dzMzMqqqqu7u7zMzM3d3d3d3d3d3d7u7u7u7u////////////////7u7u3d3d7u7u7u7u7u7u7u7u7u7uzMzMzMzMqqqqqqqqmZmZmZmZqqqqmZmZmZmZqqqqmZmZqqqqmZmZqqqqqqqqqqqqqqqqmZmZqqqqqqqqmZmZiIiIqqqqu7u7u7u7zMzMu7u7u7u7qqqqqqqqmZmZd3d3iIiImZmZu7u7u7u7u7u7u7u7qqqqqqqqzMzMzMzMzMzMzMzMzMzM3d3dzMzMzMzMqqqqqqqqqqqqqqqqu7u7qqqqmZmZd3d3d3d3iIiIqqqqu7u7zMzMzMzMzMzMqqqqqqqqmZmZmZmZmZmZmZmZqqqqmZmZmZmZmZmZiIiImZmZu7u7u7u7zMzMzMzMzMzMzMzMzMzM3d3dzMzMqqqqqqqqqqqqiIiId3d3ZmZmd3d3qqqqu7u7qqqqmZmZd3d3ZmZmZmZmZmZmZmZmd3d3d3d3iIiImZmZqqqqqqqqu7u7qqqqqqqqqqqqzMzMu7u7u7u7u7u7qqqqqqqqmZmZiIiId3d3mZmZqqqqzMzMu7u7mZmZd3d3VVVVZmZmd3d3d3d3iIiImZmZmZmZqqqqqqqqmZmZiIiId3d3ZmZmd3d3iIiIqqqqzMzMu7u7u7u7u7u7u7u7mZmZd3d3mZmZqqqqqqqqmZmZd3d3ZmZmd3d3qqqqu7u7zMzMu7u7u7u7u7u7qqqqmZmZd3d3ZmZmiIiIqqqqzMzMzMzMqqqqmZmZiIiIZmZmZmZmZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmiIiIiIiIiIiIiIiId3d3d3d3qqqqu7u7u7u7u7u7qqqqmZmZmZmZqqqqmZmZiIiIiIiIqqqqu7u7zMzMu7u7qqqqiIiId3d3u7u7zMzM3d3dzMzMqqqqmZmZd3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiImZmZu7u73d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7t3d3bu7u7u7u7u7u7u7u7u7u7u7u6qqqru7u6qqqpmZmYiIiHd3d3d3d2ZmZnd3d3d3d5mZmZmZmbu7u8zMzMzMzN3d3d3d3d3d3bu7u7u7u7u7u8zMzO7u7u7u7v///////////+7u7u7u7u7u7v///+7u7u7u7t3d3czMzLu7u6qqqpmZmZmZmZmZmYiIiJmZmYiIiJmZmZmZmZmZmZmZmaqqqqqqqqqqqpmZmZmZmZmZmYiIiHd3d4iIiIiIiKqqqru7u7u7u8zMzLu7u6qqqpmZmYiIiIiIiHd3d4iIiHd3d5mZmaqqqszMzN3d3e7u7u7u7u7u7u7u7t3d3d3d3czMzKqqqqqqqqqqqqqqqpmZmZmZmaqqqpmZmZmZmYiIiHd3d4iIiJmZmbu7u7u7u8zMzMzMzLu7u6qqqpmZmaqqqqqqqpmZmZmZmYiIiJmZmZmZmZmZmZmZmZmZmaqqqszMzMzMzN3d3d3d3czMzMzMzKqqqru7u7u7u7u7u5mZmXd3d2ZmZnd3d5mZmaqqqqqqqpmZmXd3d2ZmZmZmZlVVVWZmZnd3d3d3d5mZmYiIiIiIiKqqqqqqqpmZmaqqqru7u8zMzMzMzMzMzLu7u6qqqpmZmYiIiIiIiHd3d4iIiKqqqszMzMzMzKqqqnd3d1VVVWZmZnd3d4iIiIiIiJmZmYiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d4iIiKqqqru7u8zMzMzMzLu7u7u7u3d3d3d3d4iIiKqqqpmZmYiIiIiIiGZmZnd3d5mZmaqqqszMzMzMzMzMzMzMzKqqqpmZmXd3d3d3d3d3d5mZmbu7u7u7u7u7u6qqqnd3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZnd3d3d3d5mZmbu7u7u7u6qqqqqqqpmZmZmZmaqqqqqqqpmZmZmZmaqqqqqqqszMzLu7u6qqqoiIiIiIiJmZmczMzN3d3bu7u6qqqpmZmXd3d2ZmZmZmZnd3d4iIiHd3d3d3d4iIiJmZmaqqqszMzN3d3e7u7u7u7u7u7v///////////////+7u7v///////////////+7u7v///////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A//8AAP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////93d3bu7u8zMzMzMzMzMzLu7u7u7u7u7u7u7u6qqqqqqqqqqqpmZmYiIiIiIiHd3d3d3d3d3d6qqqru7u8zMzN3d3d3d3d3d3d3d3aqqqpmZmZmZmZmZmbu7u8zMzO7u7v///+7u7t3d3d3d3e7u7v///+7u7t3d3czMzMzMzKqqqpmZmZmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiKqqqqqqqpmZmZmZmYiIiIiIiIiIiHd3d4iIiIiIiJmZmbu7u8zMzMzMzLu7u5mZmXd3d4iIiIiIiHd3d3d3d2ZmZnd3d4iIiKqqqru7u93d3d3d3d3d3czMzMzMzKqqqqqqqpmZmZmZmaqqqpmZmZmZmZmZmZmZmZmZmaqqqoiIiIiIiHd3d5mZmaqqqru7u8zMzMzMzMzMzKqqqqqqqqqqqqqqqqqqqpmZmYiIiJmZmaqqqpmZmZmZmZmZmaqqqru7u8zMzMzMzMzMzLu7u8zMzLu7u7u7u7u7u6qqqoiIiHd3d2ZmZmZmZoiIiJmZmaqqqpmZmYiIiHd3d3d3d2ZmZmZmZmZmZnd3d4iIiIiIiJmZmZmZmZmZmaqqqqqqqru7u8zMzMzMzLu7u7u7u6qqqpmZmYiIiHd3d3d3d4iIiJmZmczMzMzMzKqqqoiIiFVVVWZmZmZmZnd3d4iIiIiIiIiIiIiIiIiIiIiIiJmZmYiIiHd3d4iIiJmZmZmZmbu7u8zMzLu7u6qqqpmZmYiIiHd3d3d3d5mZmYiIiIiIiIiIiGZmZmZmZnd3d5mZmbu7u8zMzMzMzMzMzLu7u5mZmYiIiHd3d3d3d5mZmbu7u8zMzLu7u6qqqoiIiHd3d2ZmZnd3d2ZmZlVVVWZmZmZmZnd3d3d3d3d3d4iIiHd3d3d3d2ZmZmZmZnd3d3d3d3d3d3d3d5mZmbu7u7u7u6qqqpmZmZmZmZmZmZmZmaqqqpmZmYiIiJmZmZmZmaqqqru7u6qqqoiIiIiIiJmZmczMzMzMzMzMzLu7u4iIiHd3d1VVVWZmZmZmZoiIiHd3d2ZmZmZmZoiIiKqqqru7u8zMzN3d3d3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////d3d3d3d3MzMzMzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7uqqqqZmZmZmZmZmZmZmZmZmZmZmZmqqqrMzMzd3d3d3d3MzMy7u7uqqqqIiIh3d3eIiIiZmZnMzMzd3d3d3d3d3d3d3d3u7u7u7u7d3d3d3d27u7uqqqqZmZmZmZmIiIiIiIiIiIiIiIiZmZmZmZmZmZmIiIiZmZmZmZmZmZmZmZmIiIiIiIiZmZmZmZmIiIh3d3eIiIiIiIiZmZmqqqrMzMzMzMyqqqqZmZmIiIh3d3d3d3eIiIh3d3d3d3dmZmZ3d3d3d3d3d3eIiIiZmZmqqqqqqqq7u7uqqqqZmZmqqqqqqqqZmZmIiIiIiIiIiIiZmZmqqqqZmZmIiIh3d3d3d3d3d3eZmZmqqqq7u7vMzMy7u7u7u7uqqqq7u7u7u7uqqqqqqqqZmZmZmZmqqqqqqqqqqqqZmZmZmZm7u7vMzMzMzMy7u7u7u7uqqqqqqqqqqqqqqqqZmZmZmZmIiIhmZmZmZmZmZmaZmZmqqqqqqqqZmZmZmZmIiIh3d3dmZmZ3d3d3d3d3d3eIiIiIiIiZmZmqqqqqqqqqqqqqqqq7u7u7u7u7u7u7u7uqqqqZmZmZmZl3d3d3d3d3d3eZmZm7u7u7u7u7u7uIiIh3d3dVVVVmZmZ3d3d3d3d3d3eIiIiIiIiIiIiZmZmZmZmZmZmZmZmIiIiZmZmZmZm7u7u7u7u7u7u7u7uqqqqZmZl3d3d3d3eIiIiZmZmIiIiIiIh3d3dmZmZ3d3eIiIiqqqq7u7vMzMzMzMy7u7u7u7uZmZmIiIh3d3eIiIiqqqrMzMy7u7uqqqqqqqp3d3d3d3dmZmZ3d3dmZmZmZmZ3d3d3d3eZmZmIiIh3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3eZmZmqqqqqqqqqqqqZmZl3d3d3d3eIiIiZmZmIiIiIiIiIiIiZmZmqqqqqqqqZmZmIiIh3d3eZmZm7u7vd3d3MzMyqqqqZmZl3d3dmZmZmZmZmZmZ3d3d3d3dmZmZ3d3eIiIiIiIiqqqq7u7vMzMzu7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////7u7u3d3dzMzMzMzM3d3d3d3dzMzMzMzMu7u7zMzMu7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqzMzMzMzMzMzMu7u7mZmZmZmZiIiIiIiImZmZqqqqu7u7mZmZu7u7zMzM3d3d3d3d3d3dzMzMqqqqmZmZiIiIiIiImZmZiIiImZmZmZmZmZmZmZmZmZmZmZmZmZmZiIiImZmZmZmZmZmZmZmZmZmZmZmZiIiIiIiIiIiIiIiImZmZu7u7u7u7zMzMu7u7qqqqiIiId3d3ZmZmd3d3d3d3d3d3d3d3ZmZmZmZmVVVVZmZmd3d3iIiImZmZmZmZmZmZmZmZmZmZqqqqmZmZmZmZmZmZmZmZmZmZiIiIiIiImZmZiIiId3d3iIiIiIiIqqqqu7u7u7u7u7u7qqqqqqqqqqqqzMzMu7u7qqqqmZmZmZmZmZmZqqqqmZmZqqqqmZmZu7u7u7u7u7u7qqqqu7u7qqqqqqqqmZmZmZmZmZmZqqqqiIiIZmZmZmZmd3d3mZmZu7u7u7u7qqqqiIiId3d3ZmZmd3d3d3d3iIiIiIiIiIiIiIiIiIiImZmZqqqqqqqqqqqqu7u7u7u7u7u7u7u7u7u7mZmZiIiId3d3ZmZmd3d3iIiIu7u7u7u7qqqqmZmZZmZmVVVVZmZmZmZmZmZmd3d3d3d3iIiId3d3iIiImZmZmZmZiIiImZmZmZmZqqqqqqqqu7u7zMzMqqqqqqqqiIiId3d3d3d3iIiIiIiIiIiIiIiIiIiId3d3d3d3iIiIiIiIu7u7u7u7zMzMzMzMu7u7mZmZiIiId3d3iIiIqqqqu7u7u7u7u7u7mZmZiIiIZmZmd3d3ZmZmd3d3ZmZmd3d3iIiImZmZiIiIiIiId3d3iIiImZmZiIiId3d3ZmZmZmZmZmZmmZmZqqqqu7u7mZmZd3d3ZmZmZmZmd3d3iIiId3d3iIiIiIiImZmZmZmZqqqqqqqqiIiIiIiImZmZqqqqzMzM3d3du7u7mZmZd3d3ZmZmZmZmd3d3iIiIiIiIiIiId3d3iIiImZmZqqqqu7u7zMzM7u7u////////////////////7u7u////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7t3d3czMzMzMzMzMzLu7u8zMzMzMzLu7u8zMzLu7u8zMzMzMzMzMzLu7u7u7u5mZmZmZmZmZmaqqqru7u7u7u7u7u7u7u5mZmXd3d3d3d5mZmZmZmXd3d4iIiKqqqszMzLu7u7u7u6qqqpmZmaqqqqqqqqqqqqqqqqqqqru7u6qqqqqqqpmZmaqqqpmZmZmZmZmZmZmZmZmZmZmZmaqqqpmZmZmZmZmZmYiIiJmZmZmZmYiIiIiIiJmZmbu7u93d3czMzLu7u5mZmYiIiHd3d2ZmZmZmZnd3d3d3d3d3d2ZmZmZmZlVVVWZmZnd3d3d3d4iIiIiIiIiIiJmZmYiIiJmZmaqqqpmZmYiIiJmZmYiIiJmZmYiIiHd3d3d3d3d3d4iIiJmZmbu7u7u7u7u7u6qqqqqqqqqqqru7u7u7u7u7u6qqqoiIiIiIiJmZmZmZmZmZmYiIiJmZmZmZmaqqqqqqqqqqqqqqqqqqqqqqqqqqqpmZmZmZmZmZmXd3d2ZmZnd3d6qqqru7u7u7u5mZmYiIiHd3d2ZmZnd3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiJmZmaqqqqqqqru7u7u7u7u7u7u7u7u7u5mZmYiIiHd3d3d3d3d3d3d3d5mZmbu7u7u7u6qqqnd3d1VVVVVVVVVVVVVVVWZmZnd3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiJmZmaqqqru7u8zMzLu7u6qqqpmZmXd3d2ZmZnd3d4iIiIiIiJmZmYiIiIiIiIiIiHd3d4iIiKqqqru7u8zMzMzMzLu7u6qqqoiIiHd3d3d3d5mZmbu7u7u7u7u7u6qqqoiIiGZmZnd3d3d3d3d3d2ZmZnd3d3d3d4iIiIiIiJmZmZmZmaqqqpmZmZmZmXd3d3d3d2ZmZmZmZoiIiIiIiJmZmXd3d3d3d2ZmZmZmZmZmZmZmZnd3d4iIiIiIiKqqqqqqqqqqqqqqqpmZmYiIiIiIiKqqqszMzN3d3bu7u6qqqpmZmXd3d2ZmZnd3d4iIiJmZmZmZmYiIiIiIiJmZmaqqqru7u8zMzO7u7v///////+7u7u7u7t3d3czMzMzMzO7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7d3d3MzMy7u7u7u7u7u7u7u7vMzMzMzMzMzMzMzMzd3d3d3d3MzMzMzMyqqqqIiIiIiIiZmZmqqqq7u7u7u7uqqqqIiIh3d3eIiIiZmZmqqqqIiIiZmZmqqqqZmZmZmZmZmZmZmZmZmZmqqqqqqqqqqqqqqqq7u7vMzMy7u7u7u7u7u7uqqqq7u7vMzMy7u7uqqqqqqqqqqqqZmZmZmZmZmZmZmZmZmZmqqqqZmZmIiIh3d3eZmZmqqqrMzMzd3d3d3d27u7uIiIh3d3dmZmZmZmZmZmZ3d3d3d3d3d3dmZmZ3d3dmZmZmZmZ3d3d3d3eIiIiIiIiIiIiZmZmZmZmZmZmqqqqZmZmZmZmZmZmZmZmZmZmIiIiIiIh3d3eIiIiZmZmqqqq7u7u7u7uqqqqZmZmZmZmqqqqqqqqqqqqZmZl3d3d3d3eIiIiIiIiIiIh3d3d3d3d3d3eIiIiIiIiZmZmqqqqqqqqqqqqqqqqqqqqqqqqZmZl3d3d3d3eIiIiZmZmqqqqqqqqqqqqZmZmIiIiIiIh3d3eIiIiIiIiIiIh3d3eIiIhmZmZ3d3eIiIiIiIiIiIiqqqrMzMy7u7u7u7uqqqqqqqqZmZmIiIh3d3dmZmZ3d3eZmZmqqqq7u7uqqqqIiIhVVVVEREQzMzNERERVVVVmZmZ3d3d3d3dmZmZ3d3eIiIiZmZmIiIh3d3eIiIiqqqq7u7vd3d3d3d27u7uZmZl3d3dmZmZmZmZ3d3eIiIh3d3eIiIiIiIiZmZmIiIiIiIiZmZm7u7u7u7vMzMy7u7uqqqqZmZl3d3d3d3eIiIi7u7u7u7u7u7uqqqqIiIhmZmZ3d3d3d3d3d3d3d3d3d3eIiIh3d3eZmZmqqqq7u7uqqqqZmZmZmZmIiIh3d3d3d3dVVVVmZmZ3d3eZmZmIiIh3d3dmZmZVVVVVVVVmZmZmZmZ3d3eZmZmqqqq7u7u7u7uqqqqqqqqIiIiIiIiZmZm7u7vd3d3MzMyqqqqZmZmIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3eZmZmZmZmqqqrMzMzu7u7////u7u67u7uqqqqZmZmZmZm7u7vu7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////7u7u3d3dzMzMu7u7zMzMzMzMu7u7zMzM3d3d3d3d7u7u3d3d3d3du7u7mZmZd3d3d3d3d3d3mZmZqqqqmZmZmZmZiIiIiIiImZmZqqqqu7u7qqqqmZmZiIiIiIiIiIiImZmZmZmZqqqqmZmZqqqqu7u7u7u7zMzMzMzMzMzMzMzM3d3d3d3dzMzMzMzMzMzMu7u7u7u7u7u7u7u7qqqqqqqqmZmZqqqqmZmZmZmZiIiId3d3d3d3mZmZu7u7zMzMzMzMu7u7iIiId3d3ZmZmZmZmZmZmd3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3iIiImZmZmZmZmZmZqqqqqqqqqqqqqqqqqqqqqqqqqqqqmZmZiIiIiIiId3d3iIiIiIiIqqqqu7u7zMzMu7u7qqqqmZmZiIiIiIiIiIiIiIiId3d3iIiId3d3d3d3iIiIZmZmZmZmZmZmZmZmd3d3iIiImZmZqqqqqqqqqqqqqqqqqqqqmZmZd3d3d3d3d3d3iIiImZmZqqqqqqqqqqqqmZmZiIiId3d3iIiIiIiIiIiId3d3ZmZmZmZmZmZmd3d3d3d3d3d3mZmZqqqqqqqqqqqqqqqqmZmZmZmZiIiId3d3d3d3d3d3iIiIqqqqu7u7qqqqmZmZZmZmREREMzMzMzMzREREVVVVVVVVZmZmd3d3d3d3iIiId3d3iIiId3d3iIiImZmZu7u73d3d3d3du7u7mZmZd3d3VVVVd3d3ZmZmd3d3d3d3iIiIiIiImZmZmZmZiIiImZmZqqqqu7u7zMzMzMzMu7u7iIiId3d3d3d3d3d3qqqqu7u7qqqqmZmZiIiId3d3d3d3iIiId3d3iIiId3d3iIiIiIiImZmZqqqqqqqqqqqqqqqqqqqqmZmZd3d3ZmZmZmZmZmZmiIiImZmZiIiIZmZmZmZmVVVVZmZmZmZmZmZmd3d3iIiIqqqqzMzMzMzMu7u7qqqqmZmZmZmZmZmZu7u7zMzMzMzMu7u7mZmZmZmZqqqqmZmZmZmZiIiIiIiIiIiId3d3d3d3iIiIqqqqzMzM7u7u7u7uu7u7qqqqqqqqqqqqqqqq3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////+7u7u7u7t3d3bu7u8zMzLu7u93d3d3d3e7u7t3d3d3d3czMzKqqqoiIiHd3d3d3d3d3d3d3d5mZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmYiIiHd3d3d3d3d3d4iIiJmZmaqqqqqqqru7u7u7u7u7u8zMzMzMzMzMzN3d3d3d3d3d3czMzN3d3czMzMzMzMzMzMzMzMzMzMzMzLu7u6qqqpmZmZmZmaqqqpmZmXd3d3d3d3d3d5mZmaqqqszMzLu7u4iIiGZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiIiIiIiIiJmZmYiIiJmZmaqqqqqqqru7u6qqqqqqqqqqqru7u6qqqqqqqqqqqpmZmZmZmZmZmYiIiHd3d4iIiKqqqru7u8zMzLu7u6qqqpmZmYiIiHd3d5mZmZmZmYiIiHd3d2ZmZlVVVWZmZmZmZmZmZlVVVVVVVVVVVYiIiJmZmaqqqru7u6qqqqqqqqqqqoiIiHd3d3d3d3d3d3d3d5mZmaqqqru7u7u7u5mZmXd3d3d3d4iIiIiIiIiIiIiIiGZmZlVVVVVVVVVVVWZmZmZmZoiIiIiIiJmZmZmZmZmZmZmZmYiIiHd3d3d3d2ZmZnd3d4iIiKqqqru7u7u7u5mZmWZmZkRERCIiIjMzMzMzM0RERFVVVWZmZnd3d3d3d3d3d4iIiHd3d3d3d4iIiIiIiLu7u8zMzMzMzLu7u5mZmXd3d2ZmZmZmZmZmZnd3d3d3d4iIiJmZmaqqqpmZmZmZmZmZmaqqqqqqqru7u7u7u6qqqoiIiHd3d2ZmZmZmZoiIiLu7u7u7u6qqqoiIiIiIiHd3d3d3d3d3d3d3d3d3d4iIiJmZmYiIiJmZmaqqqru7u7u7u7u7u5mZmYiIiHd3d2ZmZmZmZnd3d3d3d3d3d3d3d4iIiHd3d1VVVVVVVWZmZnd3d4iIiKqqqszMzMzMzLu7u6qqqpmZmZmZmZmZmbu7u7u7u8zMzKqqqru7u7u7u8zMzLu7u4iIiIiIiIiIiIiIiHd3d2ZmZnd3d4iIiLu7u+7u7t3d3czMzMzMzLu7u7u7u7u7u93d3f///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////u7u7////////////////////u7u7////////////////////u7u7////u7u7u7u7MzMzMzMzu7u7u7u7////////////////////////////////////////////////////////////////////////////u7u7d3d3d3d3MzMzd3d3d3d3d3d3u7u7MzMy7u7uZmZmZmZl3d3dmZmZmZmZmZmZ3d3eZmZmqqqqqqqq7u7uqqqqqqqqZmZmZmZmIiIh3d3dmZmZ3d3d3d3eZmZmZmZmqqqq7u7u7u7u7u7vMzMzMzMzd3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMy7u7uqqqqqqqq7u7uZmZmIiIhmZmZ3d3eIiIiqqqq7u7uqqqqZmZmIiIiIiIh3d3dmZmZ3d3d3d3eIiIiIiIiIiIiZmZmqqqqqqqqqqqqqqqqqqqq7u7u7u7uqqqqqqqq7u7u7u7vMzMyqqqqqqqqqqqqZmZmIiIiIiIiIiIh3d3eZmZmqqqrMzMy7u7u7u7uZmZmIiIh3d3eZmZmZmZl3d3dmZmZERERVVVVVVVV3d3d3d3dmZmZVVVVVVVVmZmZ3d3eqqqqqqqqqqqqZmZmZmZmIiIiZmZl3d3dmZmZ3d3d3d3eqqqq7u7u7u7uZmZmIiIh3d3d3d3eIiIiIiIiIiIhmZmZERERERERERERVVVVVVVVmZmaIiIiZmZmZmZmZmZmIiIiIiIiIiIhmZmZmZmZmZmZ3d3eZmZm7u7u7u7uqqqp3d3dVVVUzMzMzMzMzMzNERERERERVVVVmZmZ3d3d3d3eIiIiIiIh3d3d3d3eIiIi7u7u7u7u7u7uqqqqZmZl3d3dmZmZmZmZmZmZmZmZ3d3d3d3eIiIiqqqqqqqqZmZmIiIiZmZmqqqqqqqqqqqqqqqqZmZl3d3dmZmZmZmaIiIiqqqq7u7uqqqqZmZl3d3dmZmZ3d3d3d3d3d3d3d3eIiIiZmZmZmZmZmZmqqqq7u7u7u7u7u7uqqqqIiIhmZmZmZmZmZmZmZmZ3d3eIiIiIiIhmZmZERERERERVVVVmZmZmZmZmZmaqqqrMzMzd3d3MzMy7u7uqqqqZmZmqqqqqqqq7u7vMzMzMzMzMzMzMzMzMzMy7u7uZmZmIiIiIiIh3d3dmZmZVVVVmZmaIiIi7u7vd3d3MzMzMzMy7u7u7u7uqqqrMzMzd3d3////////////////////u7u7////////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////7u7u////7u7u7u7u7u7u7u7u7u7u7u7u////////////////7u7u7u7u3d3du7u7u7u7qqqqzMzM7u7u7u7u////////////7u7u7u7u7u7u7u7u////////7u7u////7u7u////7u7u////7u7u////////////7u7u7u7u3d3d7u7u7u7u3d3d3d3du7u7qqqqmZmZiIiId3d3d3d3VVVVZmZmZmZmiIiImZmZqqqqu7u7u7u7u7u7qqqqqqqqmZmZiIiId3d3ZmZmd3d3d3d3iIiIqqqqzMzMzMzMzMzMu7u7zMzM3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d7u7u7u7u3d3d3d3dzMzMzMzMu7u7u7u7qqqqqqqqmZmZd3d3ZmZmd3d3mZmZqqqqqqqqqqqqmZmZiIiIiIiIZmZmZmZmd3d3d3d3iIiImZmZqqqqqqqqu7u7qqqqqqqqmZmZmZmZu7u7u7u7u7u7u7u7zMzMzMzMzMzMu7u7qqqqqqqqiIiIiIiId3d3d3d3iIiIqqqqu7u7u7u7u7u7mZmZmZmZd3d3iIiIiIiIiIiIVVVVVVVVREREVVVViIiImZmZiIiIZmZmVVVVZmZmd3d3mZmZqqqqmZmZiIiIiIiImZmZiIiId3d3ZmZmd3d3iIiIqqqqu7u7qqqqiIiIiIiId3d3d3d3d3d3mZmZiIiIZmZmVVVVMzMzMzMzREREREREZmZmd3d3d3d3mZmZmZmZmZmZiIiId3d3ZmZmVVVVZmZmd3d3iIiIqqqqzMzMu7u7mZmZZmZmMzMzMzMzMzMzREREMzMzVVVVVVVVZmZmZmZmd3d3d3d3iIiId3d3iIiImZmZu7u7u7u7qqqqiIiIZmZmVVVVVVVVZmZmd3d3d3d3d3d3iIiImZmZmZmZiIiIiIiIiIiImZmZmZmZqqqqmZmZmZmZd3d3ZmZmZmZmd3d3mZmZqqqqqqqqiIiIiIiId3d3ZmZmZmZmd3d3d3d3iIiIiIiIiIiImZmZiIiIqqqqzMzMzMzMu7u7mZmZd3d3ZmZmZmZmZmZmd3d3iIiId3d3VVVVREREVVVVVVVVVVVVVVVVZmZmmZmZzMzM3d3d3d3du7u7qqqqmZmZmZmZu7u7u7u7zMzMzMzMu7u7u7u7zMzMzMzMqqqqiIiIiIiId3d3ZmZmZmZmZmZmiIiIqqqqzMzMzMzMu7u7u7u7mZmZmZmZqqqqzMzM7u7u////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7u7u7t3d3d3d3d3d3czMzMzMzLu7u6qqqqqqqru7u93d3e7u7u7u7v///////+7u7u7u7t3d3bu7u6qqqru7u7u7u8zMzO7u7u7u7v///////+7u7t3d3e7u7t3d3e7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3e7u7u7u7u7u7u7u7u7u7u7u7t3d3czMzKqqqpmZmYiIiIiIiJmZmXd3d3d3d2ZmZnd3d3d3d5mZmbu7u7u7u8zMzLu7u7u7u6qqqpmZmYiIiHd3d3d3d3d3d3d3d5mZmaqqqru7u7u7u7u7u8zMzMzMzMzMzN3d3czMzN3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzLu7u7u7u7u7u6qqqoiIiHd3d2ZmZnd3d4iIiKqqqqqqqpmZmZmZmYiIiHd3d3d3d2ZmZnd3d3d3d4iIiIiIiJmZmbu7u7u7u7u7u6qqqpmZmZmZmbu7u7u7u7u7u8zMzMzMzMzMzMzMzLu7u7u7u6qqqpmZmZmZmXd3d3d3d4iIiJmZmbu7u8zMzLu7u6qqqpmZmXd3d3d3d4iIiHd3d2ZmZlVVVVVVVXd3d5mZmaqqqpmZmXd3d3d3d3d3d4iIiJmZmZmZmYiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d4iIiJmZmaqqqqqqqpmZmYiIiHd3d3d3d3d3d3d3d3d3d3d3d1VVVTMzMzMzMzMzM0RERERERFVVVWZmZoiIiJmZmZmZmYiIiIiIiGZmZmZmZlVVVWZmZoiIiKqqqru7u7u7u5mZmWZmZlVVVTMzMzMzM0RERDMzM0RERFVVVWZmZnd3d3d3d4iIiIiIiHd3d4iIiJmZmbu7u7u7u5mZmXd3d3d3d2ZmZlVVVWZmZmZmZmZmZmZmZnd3d4iIiIiIiJmZmYiIiHd3d4iIiJmZmZmZmYiIiHd3d3d3d2ZmZmZmZmZmZoiIiKqqqqqqqqqqqpmZmXd3d3d3d3d3d3d3d3d3d3d3d4iIiJmZmYiIiJmZmaqqqru7u8zMzLu7u5mZmYiIiGZmZmZmZnd3d3d3d4iIiHd3d1VVVVVVVVVVVURERERERFVVVWZmZpmZmbu7u93d3czMzMzMzKqqqpmZmZmZmaqqqszMzMzMzMzMzLu7u7u7u7u7u7u7u6qqqoiIiHd3d3d3d3d3d3d3d3d3d4iIiKqqqru7u7u7u6qqqqqqqpmZmZmZmZmZmczMzO7u7v///+7u7u7u7v///+7u7v///////////+7u7v///////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////u7u7////u7u7u7u7d3d3d3d3MzMzMzMy7u7uqqqqZmZmZmZmZmZmZmZmqqqq7u7vMzMzd3d3d3d3////u7u7////u7u7MzMzMzMyqqqqqqqq7u7u7u7vMzMzu7u7////u7u7u7u7u7u7d3d3d3d3u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7////u7u7u7u7d3d27u7uqqqqZmZmZmZmqqqqZmZmZmZl3d3d3d3d3d3eIiIiZmZm7u7u7u7vMzMzMzMzMzMy7u7uqqqqZmZmZmZmIiIiIiIh3d3eIiIiZmZmqqqq7u7u7u7u7u7u7u7vMzMzd3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3d3d3d3d3d3d3MzMzMzMzMzMy7u7uqqqqqqqqZmZmIiIh3d3dmZmZ3d3eZmZm7u7uqqqqZmZmIiIh3d3dmZmZmZmZmZmZ3d3eIiIiIiIiqqqqqqqq7u7u7u7u7u7uqqqqqqqq7u7u7u7vMzMzd3d3MzMzMzMy7u7vMzMzMzMy7u7uqqqqZmZl3d3eIiIiIiIiZmZmqqqrMzMy7u7u7u7uZmZmIiIh3d3d3d3d3d3dmZmZVVVVVVVVmZmaIiIiqqqqIiIiZmZmIiIiIiIiIiIiIiIh3d3d3d3eIiIiIiIiZmZmZmZmIiIh3d3d3d3eIiIiZmZmqqqqqqqqqqqqZmZl3d3d3d3d3d3eIiIiIiIiIiIhmZmZEREQzMzMiIiIzMzMzMzNERERVVVWIiIiIiIiIiIiIiIiIiIhmZmZmZmZVVVVmZmaIiIiqqqq7u7u7u7uqqqqIiIhmZmZEREQzMzMzMzMzMzNERERERERVVVV3d3eZmZmZmZmIiIiIiIiIiIiZmZmqqqq7u7u7u7uZmZl3d3dVVVVVVVVmZmZmZmZ3d3d3d3dmZmZ3d3eZmZmZmZmZmZmIiIh3d3eIiIiIiIh3d3dmZmZmZmZmZmZVVVVmZmaIiIiqqqq7u7uqqqqZmZl3d3eIiIiIiIh3d3d3d3d3d3eIiIiZmZmZmZmqqqqqqqq7u7vMzMyqqqqqqqqIiIhmZmZmZmZ3d3eIiIiIiIh3d3dmZmZERERERERVVVVERERVVVVmZmaIiIiZmZnMzMzMzMy7u7uqqqqZmZmZmZmqqqrMzMzMzMy7u7vMzMyqqqq7u7uqqqqqqqqIiIh3d3dmZmZ3d3eIiIiIiIiIiIiZmZmqqqqqqqqqqqqZmZmZmZmIiIiZmZm7u7vd3d3u7u7d3d3d3d3MzMzd3d3u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3dzMzMu7u7u7u7qqqqqqqqqqqqmZmZqqqqqqqqu7u7zMzM3d3d7u7u7u7u////3d3d3d3dzMzMu7u7u7u7u7u7u7u7zMzM3d3d3d3d7u7u7u7u3d3d3d3d3d3d7u7u7u7u////////7u7u////7u7u7u7u7u7u7u7u////7u7u7u7u7u7u7u7u3d3dzMzMu7u7u7u7u7u7qqqqqqqqmZmZiIiIiIiId3d3iIiIiIiImZmZu7u7zMzMzMzMzMzMu7u7qqqqqqqqqqqqmZmZmZmZiIiIiIiId3d3mZmZqqqqu7u7u7u7u7u7zMzMzMzMzMzMzMzMzMzM3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3dzMzMzMzMu7u7u7u7qqqqqqqqmZmZd3d3ZmZmd3d3mZmZqqqqu7u7qqqqiIiId3d3ZmZmZmZmZmZmd3d3d3d3iIiImZmZmZmZqqqqu7u7zMzMu7u7u7u7u7u7u7u7zMzM3d3d3d3d3d3dzMzMzMzM3d3d3d3du7u7qqqqiIiIiIiId3d3iIiImZmZu7u7zMzMu7u7qqqqiIiId3d3d3d3iIiId3d3ZmZmREREVVVVd3d3iIiId3d3iIiImZmZiIiIiIiId3d3ZmZmd3d3iIiIiIiImZmZmZmZmZmZiIiIiIiIiIiImZmZmZmZqqqqmZmZmZmZiIiId3d3d3d3iIiImZmZiIiId3d3VVVVMzMzREREREREMzMzREREVVVVZmZmd3d3d3d3iIiId3d3d3d3ZmZmVVVVZmZmZmZmmZmZu7u7u7u7u7u7mZmZd3d3ZmZmREREREREREREREREVVVVZmZmd3d3mZmZmZmZmZmZiIiId3d3iIiIqqqqu7u7u7u7mZmZiIiIZmZmVVVVVVVVd3d3d3d3d3d3ZmZmZmZmiIiImZmZiIiIiIiIiIiIiIiId3d3iIiId3d3ZmZmZmZmVVVVVVVVd3d3mZmZqqqqu7u7qqqqmZmZiIiIiIiId3d3iIiId3d3ZmZmiIiImZmZqqqqqqqqu7u7zMzMu7u7qqqqmZmZd3d3ZmZmd3d3d3d3iIiId3d3VVVVVVVVREREREREVVVVVVVVZmZmZmZmiIiIqqqqzMzMu7u7qqqqmZmZqqqqqqqqu7u7u7u7zMzMzMzMu7u7qqqqqqqqmZmZiIiId3d3ZmZmd3d3mZmZiIiIiIiImZmZiIiImZmZmZmZmZmZmZmZmZmZiIiIqqqqzMzM3d3dzMzMu7u7qqqqu7u73d3d////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7t3d3e7u7u7u7u7u7t3d3d3d3d3d3e7u7u7u7u7u7u7u7t3d3e7u7t3d3czMzMzMzLu7u7u7u6qqqqqqqqqqqru7u7u7u93d3d3d3d3d3e7u7t3d3d3d3czMzMzMzLu7u7u7u7u7u7u7u7u7u8zMzMzMzLu7u7u7u93d3e7u7u7u7u7u7v///+7u7v///////////////////+7u7u7u7t3d3d3d3d3d3d3d3czMzMzMzMzMzLu7u7u7u6qqqqqqqqqqqpmZmXd3d3d3d3d3d5mZmaqqqru7u8zMzLu7u8zMzLu7u6qqqqqqqqqqqpmZmYiIiIiIiIiIiJmZmaqqqru7u6qqqru7u8zMzMzMzMzMzMzMzN3d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3czMzLu7u7u7u7u7u7u7u6qqqpmZmXd3d2ZmZnd3d4iIiJmZmaqqqru7u5mZmYiIiGZmZmZmZmZmZnd3d4iIiHd3d4iIiIiIiJmZmbu7u8zMzMzMzLu7u7u7u7u7u8zMzN3d3d3d3czMzN3d3d3d3d3d3czMzLu7u5mZmYiIiHd3d3d3d3d3d5mZmbu7u8zMzLu7u6qqqoiIiIiIiHd3d3d3d4iIiGZmZlVVVVVVVWZmZnd3d3d3d3d3d5mZmYiIiIiIiIiIiIiIiIiIiHd3d4iIiIiIiKqqqqqqqqqqqoiIiJmZmYiIiJmZmZmZmZmZmYiIiHd3d3d3d3d3d5mZmZmZmYiIiHd3d1VVVVVVVVVVVURERERERERERERERFVVVWZmZnd3d4iIiIiIiHd3d2ZmZlVVVVVVVWZmZpmZmbu7u7u7u7u7u5mZmXd3d2ZmZlVVVWZmZlVVVURERFVVVXd3d3d3d5mZmZmZmZmZmYiIiIiIiIiIiKqqqru7u7u7u6qqqnd3d1VVVVVVVVVVVXd3d4iIiHd3d2ZmZlVVVWZmZoiIiJmZmYiIiHd3d3d3d3d3d3d3d3d3d2ZmZmZmZlVVVVVVVWZmZoiIiLu7u7u7u6qqqpmZmYiIiHd3d4iIiIiIiHd3d3d3d3d3d5mZmZmZmaqqqru7u8zMzLu7u6qqqoiIiHd3d2ZmZmZmZmZmZoiIiHd3d1VVVVVVVVVVVURERFVVVXd3d2ZmZnd3d4iIiKqqqru7u8zMzKqqqqqqqpmZmaqqqszMzMzMzMzMzLu7u6qqqqqqqqqqqqqqqpmZmXd3d3d3d4iIiKqqqqqqqpmZmYiIiIiIiJmZmaqqqpmZmZmZmZmZmYiIiKqqqru7u6qqqqqqqqqqqru7u6qqqt3d3e7u7v///////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////d3d3d3d3d3d3u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3MzMzMzMzMzMy7u7uqqqqqqqqqqqqqqqq7u7u7u7u7u7vd3d3d3d3u7u7d3d3MzMy7u7u7u7uqqqqIiIiZmZmZmZmIiIiZmZnMzMzd3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7////u7u7////u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMy7u7vMzMy7u7u7u7uZmZmIiIiIiIiIiIiIiIiZmZmqqqq7u7u7u7u7u7u7u7u7u7uqqqqZmZmZmZmZmZmZmZmIiIiZmZmZmZmqqqq7u7vMzMy7u7vMzMy7u7vMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMy7u7u7u7u7u7uqqqqqqqqZmZmIiIhmZmZmZmZ3d3eZmZmqqqq7u7uqqqqIiIiIiIh3d3dmZmZmZmZ3d3eIiIiIiIiIiIiIiIiZmZm7u7vMzMzMzMy7u7vMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyqqqqqqqqIiIh3d3d3d3d3d3eIiIiqqqq7u7u7u7u7u7uZmZmIiIhmZmZ3d3eIiIh3d3dmZmZVVVVmZmZ3d3eIiIiIiIiZmZmqqqqqqqqqqqqZmZmZmZmZmZmZmZm7u7uqqqq7u7uqqqqZmZmIiIiIiIiZmZmZmZmIiIh3d3d3d3dmZmaIiIiIiIiIiIiZmZl3d3dmZmZVVVVVVVVVVVVmZmZVVVVERERVVVVVVVWIiIiIiIh3d3d3d3dmZmZVVVVVVVVmZmZ3d3eqqqq7u7uqqqqZmZl3d3dmZmZ3d3eIiIh3d3dVVVVVVVVmZmaIiIiIiIiZmZmqqqqZmZl3d3eIiIiZmZmqqqrMzMyqqqp3d3dmZmZVVVVmZmZ3d3eIiIiIiIhmZmZERERmZmZ3d3d3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3dmZmZVVVVVVVVmZmaIiIiqqqq7u7u7u7uZmZmIiIh3d3eIiIiZmZmIiIh3d3d3d3d3d3eZmZm7u7vMzMy7u7uqqqqZmZmIiIhmZmZmZmZVVVV3d3eZmZl3d3dmZmZVVVVVVVVmZmZ3d3d3d3dmZmZmZmaIiIiqqqq7u7vMzMy7u7uqqqqZmZm7u7u7u7vMzMy7u7u7u7uZmZmZmZmqqqq7u7uqqqqIiIh3d3eZmZm7u7u7u7uZmZmZmZmZmZmZmZmZmZmqqqqqqqqqqqqZmZmIiIiIiIiIiIiZmZmZmZmZmZmqqqrMzMzu7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3d3d3d7u7u7u7u3d3d7u7u7u7u////7u7u////7u7u7u7u7u7u7u7u3d3dzMzMzMzMzMzMzMzMzMzMu7u7qqqqqqqqmZmZmZmZiIiImZmZiIiImZmZqqqqzMzM3d3d3d3d3d3dzMzMzMzMu7u7qqqqiIiId3d3d3d3mZmZmZmZu7u7u7u7u7u7u7u7zMzM3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3dzMzM3d3d7u7u7u7u3d3d3d3dzMzMzMzMu7u7u7u7mZmZiIiId3d3d3d3d3d3iIiImZmZqqqqu7u7zMzMzMzMu7u7u7u7qqqqmZmZmZmZmZmZmZmZiIiIiIiImZmZu7u7u7u7u7u7u7u7zMzMzMzMu7u7zMzMzMzMzMzM3d3d3d3d3d3dzMzMzMzMu7u7u7u7u7u7qqqqqqqqqqqqmZmZiIiId3d3d3d3d3d3iIiImZmZqqqqqqqqmZmZiIiId3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiIqqqqu7u7zMzMzMzM3d3dzMzMzMzMu7u7zMzMzMzMzMzMzMzMu7u7u7u7qqqqmZmZd3d3d3d3ZmZmiIiIiIiIu7u7u7u7u7u7qqqqd3d3ZmZmZmZmd3d3d3d3d3d3ZmZmZmZmiIiIiIiIqqqqu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7qqqqqqqqmZmZiIiIiIiIiIiIiIiImZmZiIiId3d3ZmZmd3d3iIiIiIiIiIiId3d3ZmZmVVVVZmZmd3d3d3d3ZmZmVVVVVVVVVVVVZmZmd3d3iIiIiIiIZmZmZmZmVVVVVVVVd3d3mZmZu7u7u7u7qqqqiIiId3d3iIiIiIiIiIiId3d3ZmZmVVVVd3d3iIiImZmZmZmZmZmZiIiIiIiImZmZqqqqzMzMu7u7mZmZd3d3ZmZmd3d3ZmZmiIiId3d3d3d3ZmZmVVVVZmZmZmZmd3d3iIiId3d3d3d3d3d3iIiId3d3VVVVVVVVVVVVVVVVd3d3mZmZu7u7u7u7mZmZd3d3d3d3d3d3iIiIiIiIZmZmZmZmZmZmmZmZqqqqu7u7qqqqmZmZmZmZd3d3ZmZmVVVVZmZmd3d3iIiIiIiId3d3VVVVZmZmd3d3ZmZmd3d3d3d3d3d3d3d3mZmZqqqqu7u7u7u7qqqqqqqqqqqqu7u7u7u7u7u7u7u7qqqqmZmZmZmZu7u7qqqqmZmZiIiImZmZqqqqu7u7qqqqqqqqmZmZmZmZmZmZu7u7zMzMqqqqmZmZiIiId3d3d3d3d3d3iIiIiIiImZmZu7u7zMzM7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7u7u7u7u7v///+7u7u7u7u7u7t3d3d3d3bu7u7u7u7u7u6qqqru7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqqqqqpmZmZmZmYiIiIiIiHd3d4iIiKqqqru7u93d3d3d3czMzN3d3czMzLu7u5mZmYiIiIiIiIiIiIiIiIiIiIiIiJmZmaqqqszMzMzMzMzMzMzMzN3d3czMzN3d3czMzN3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzLu7u5mZmZmZmYiIiHd3d3d3d2ZmZnd3d4iIiJmZmaqqqru7u7u7u8zMzLu7u6qqqqqqqpmZmZmZmZmZmZmZmZmZmaqqqpmZmZmZmaqqqru7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u8zMzN3d3bu7u7u7u6qqqqqqqqqqqqqqqpmZmZmZmYiIiHd3d3d3d2ZmZnd3d4iIiJmZmaqqqoiIiIiIiHd3d4iIiIiIiIiIiIiIiHd3d3d3d3d3d4iIiJmZmaqqqru7u8zMzMzMzMzMzN3d3czMzMzMzLu7u7u7u7u7u7u7u6qqqpmZmYiIiHd3d3d3d2ZmZnd3d4iIiKqqqru7u7u7u6qqqnd3d3d3d3d3d3d3d4iIiHd3d3d3d2ZmZnd3d5mZmbu7u7u7u8zMzLu7u8zMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u6qqqpmZmYiIiIiIiIiIiIiIiIiIiIiIiGZmZmZmZmZmZnd3d4iIiIiIiIiIiGZmZmZmZmZmZnd3d3d3d4iIiHd3d1VVVURERERERGZmZnd3d3d3d3d3d1VVVVVVVWZmZnd3d5mZmaqqqru7u7u7u5mZmYiIiIiIiKqqqqqqqpmZmXd3d2ZmZmZmZmZmZnd3d5mZmZmZmYiIiIiIiIiIiJmZmbu7u8zMzKqqqoiIiIiIiHd3d3d3d4iIiIiIiHd3d2ZmZlVVVVVVVWZmZmZmZmZmZnd3d3d3d4iIiHd3d2ZmZlVVVWZmZlVVVVVVVWZmZpmZmaqqqqqqqpmZmXd3d2ZmZnd3d4iIiIiIiGZmZmZmZlVVVVVVVXd3d5mZmaqqqqqqqoiIiGZmZmZmZlVVVWZmZnd3d4iIiIiIiHd3d2ZmZmZmZmZmZmZmZmZmZoiIiHd3d3d3d5mZmZmZmaqqqru7u7u7u5mZmaqqqqqqqru7u8zMzLu7u6qqqqqqqqqqqru7u6qqqpmZmYiIiJmZmaqqqszMzLu7u6qqqpmZmYiIiJmZmczMzMzMzLu7u5mZmYiIiHd3d3d3d4iIiHd3d2ZmZoiIiJmZmczMzN3d3e7u7v///+7u7v///////+7u7v///////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7////u7u7u7u7u7u7u7u7MzMy7u7uZmZmZmZmZmZmqqqqqqqqqqqqqqqqqqqqqqqq7u7u7u7vMzMzMzMzMzMyqqqqZmZmZmZmIiIh3d3eIiIiIiIi7u7vMzMzd3d3d3d3MzMzMzMyqqqqZmZmIiIh3d3d3d3dmZmZ3d3d3d3eIiIiZmZmqqqq7u7u7u7u7u7vMzMy7u7vMzMzMzMy7u7vMzMzMzMzMzMzMzMzd3d3d3d3MzMzMzMzMzMzMzMyqqqqqqqqZmZmIiIh3d3d3d3d3d3d3d3d3d3d3d3eIiIiZmZmqqqq7u7u7u7u7u7u7u7uqqqqZmZmZmZmqqqqZmZmqqqqZmZmZmZmIiIiqqqqqqqq7u7u7u7u7u7uqqqqqqqqZmZmZmZmqqqq7u7vMzMy7u7uqqqqqqqqqqqqZmZmZmZmqqqqqqqqIiIh3d3d3d3dmZmZ3d3eZmZmZmZmZmZmZmZl3d3d3d3d3d3eIiIh3d3dmZmZ3d3eIiIiIiIiIiIiZmZmqqqq7u7vMzMzd3d3MzMzd3d3d3d3d3d3MzMy7u7uqqqqqqqqZmZmIiIiIiIh3d3d3d3d3d3d3d3eIiIiZmZmZmZmqqqqqqqqqqqqZmZl3d3dmZmaIiIh3d3eIiIh3d3eIiIiZmZmqqqq7u7vMzMzMzMzMzMy7u7vMzMzMzMzMzMzMzMzMzMzMzMy7u7uZmZmIiIiIiIiIiIiZmZmIiIiIiIh3d3d3d3d3d3eIiIiIiIiIiIh3d3d3d3dmZmZmZmZmZmZ3d3eIiIiIiIhmZmZVVVVVVVVmZmZ3d3d3d3dmZmZmZmZVVVVmZmZ3d3eIiIiqqqrMzMy7u7uqqqqZmZmZmZmZmZm7u7uZmZl3d3dmZmZVVVVmZmZmZmZ3d3eZmZmZmZmIiIiIiIiZmZmqqqqqqqqZmZmZmZmIiIiIiIh3d3d3d3d3d3d3d3dmZmZmZmZERERVVVVVVVV3d3d3d3eIiIiIiIh3d3dmZmZmZmZmZmZVVVVVVVVmZmaIiIiqqqqqqqqZmZmIiIh3d3dmZmZ3d3eIiIh3d3dVVVVERERVVVVmZmZ3d3eIiIiZmZl3d3dmZmZVVVVVVVVmZmZ3d3eIiIiIiIh3d3dmZmZmZmZVVVV3d3d3d3eIiIh3d3d3d3eIiIiIiIiqqqq7u7u7u7uqqqqqqqq7u7u7u7u7u7vMzMy7u7u7u7uqqqq7u7uqqqqZmZmZmZmZmZm7u7vMzMy7u7uqqqqZmZmZmZm7u7vMzMzMzMy7u7uqqqqIiIiIiIiIiIiqqqqIiIh3d3d3d3eqqqrMzMzd3d3u7u7////////////////////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u3d3du7u7qqqqmZmZqqqqqqqqqqqqmZmZmZmZiIiImZmZqqqqu7u7u7u7u7u7zMzMzMzMzMzMu7u7qqqqmZmZiIiId3d3iIiImZmZqqqqzMzM3d3dzMzMzMzMu7u7qqqqiIiId3d3ZmZmZmZmZmZmZmZmZmZmd3d3mZmZu7u7zMzMu7u7zMzMzMzMu7u7u7u7zMzM3d3dzMzM3d3dzMzMzMzMzMzMzMzMu7u7u7u7qqqqu7u7mZmZmZmZiIiIiIiId3d3d3d3d3d3d3d3ZmZmd3d3iIiIqqqqqqqqu7u7u7u7u7u7qqqqqqqqmZmZmZmZqqqqqqqqqqqqmZmZiIiImZmZiIiImZmZqqqqu7u7u7u7qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqmZmZmZmZmZmZmZmZqqqqiIiIiIiId3d3ZmZmd3d3d3d3iIiIiIiIiIiId3d3iIiIiIiIiIiIZmZmZmZmd3d3iIiIiIiId3d3d3d3mZmZqqqqu7u7zMzM3d3d3d3d3d3dzMzMzMzMu7u7qqqqmZmZiIiIiIiIZmZmZmZmd3d3d3d3d3d3d3d3iIiImZmZzMzMzMzMu7u7mZmZd3d3d3d3d3d3mZmZiIiIiIiIiIiImZmZqqqqqqqqzMzMzMzMzMzMzMzMzMzMzMzM3d3dzMzM3d3dzMzMu7u7qqqqiIiIiIiIiIiImZmZiIiIiIiId3d3ZmZmd3d3d3d3iIiImZmZiIiId3d3d3d3d3d3iIiIiIiImZmZmZmZd3d3ZmZmZmZmZmZmd3d3d3d3d3d3d3d3ZmZmd3d3d3d3iIiIqqqqzMzMu7u7u7u7mZmZiIiImZmZu7u7qqqqiIiIZmZmZmZmVVVVZmZmiIiIiIiIiIiIiIiId3d3iIiIqqqqmZmZmZmZmZmZmZmZiIiIiIiId3d3d3d3d3d3d3d3VVVVVVVVVVVVZmZmd3d3d3d3d3d3iIiIiIiId3d3ZmZmZmZmVVVVVVVVZmZmZmZmmZmZqqqqqqqqmZmZZmZmZmZmZmZmd3d3d3d3VVVVREREREREREREZmZmZmZmd3d3d3d3d3d3d3d3VVVVZmZmd3d3d3d3d3d3d3d3ZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3iIiImZmZmZmZu7u7u7u7qqqqmZmZqqqqu7u7zMzMu7u7zMzMu7u7qqqqu7u7u7u7qqqqqqqqmZmZu7u7u7u7zMzMu7u7mZmZmZmZu7u73d3dzMzMqqqqmZmZiIiIiIiImZmZqqqqmZmZiIiIiIiIqqqqu7u7zMzM7u7u7u7u////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7u7u7t3d3czMzKqqqpmZmaqqqpmZmaqqqpmZmZmZmZmZmZmZmZmZmZmZmZmZmaqqqpmZmbu7u8zMzMzMzLu7u6qqqqqqqpmZmYiIiIiIiIiIiJmZmaqqqru7u93d3d3d3czMzLu7u6qqqoiIiHd3d2ZmZmZmZmZmZmZmZnd3d4iIiJmZmaqqqru7u7u7u7u7u7u7u7u7u8zMzMzMzMzMzLu7u8zMzMzMzMzMzKqqqqqqqpmZmZmZmZmZmZmZmYiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d2ZmZnd3d4iIiJmZmbu7u7u7u7u7u7u7u5mZmYiIiJmZmZmZmaqqqpmZmZmZmYiIiHd3d3d3d4iIiJmZmZmZmaqqqqqqqpmZmZmZmZmZmZmZmYiIiIiIiIiIiIiIiJmZmZmZmZmZmaqqqpmZmYiIiIiIiIiIiHd3d3d3d2ZmZoiIiIiIiJmZmaqqqqqqqoiIiGZmZmZmZmZmZnd3d4iIiHd3d3d3d3d3d3d3d4iIiJmZmbu7u8zMzN3d3d3d3bu7u7u7u6qqqqqqqpmZmYiIiIiIiHd3d1VVVWZmZmZmZmZmZmZmZnd3d5mZmaqqqszMzKqqqpmZmXd3d4iIiIiIiJmZmZmZmZmZmZmZmZmZmZmZmaqqqru7u7u7u8zMzMzMzMzMzMzMzMzMzN3d3czMzMzMzLu7u6qqqoiIiIiIiHd3d5mZmZmZmYiIiGZmZmZmZnd3d3d3d4iIiJmZmZmZmYiIiGZmZnd3d5mZmaqqqru7u7u7u6qqqoiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d2ZmZnd3d4iIiKqqqru7u7u7u6qqqpmZmYiIiJmZmbu7u7u7u5mZmXd3d2ZmZmZmZmZmZnd3d5mZmZmZmYiIiHd3d5mZmZmZmYiIiKqqqpmZmXd3d2ZmZnd3d4iIiIiIiIiIiGZmZmZmZlVVVVVVVWZmZmZmZnd3d3d3d3d3d5mZmYiIiIiIiHd3d1VVVWZmZmZmZmZmZoiIiKqqqqqqqpmZmXd3d1VVVWZmZnd3d3d3d2ZmZkRERERERERERERERGZmZnd3d3d3d4iIiHd3d2ZmZmZmZmZmZoiIiIiIiIiIiGZmZmZmZnd3d2ZmZnd3d3d3d3d3d4iIiIiIiIiIiJmZmaqqqru7u6qqqpmZmaqqqru7u7u7u8zMzLu7u7u7u7u7u7u7u7u7u7u7u6qqqqqqqqqqqru7u8zMzKqqqoiIiJmZmbu7u8zMzKqqqqqqqqqqqpmZmYiIiIiIiKqqqqqqqoiIiIiIiKqqqru7u8zMzO7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////u7u7////////////////////////////////////////////u7u7u7u7u7u7MzMyqqqqIiIiIiIiZmZmZmZmZmZmZmZmZmZmZmZmIiIiqqqqZmZmqqqqZmZmZmZmZmZm7u7u7u7u7u7uqqqqqqqqIiIiZmZmIiIiIiIiIiIiqqqqqqqq7u7vd3d3MzMzMzMyqqqqqqqqZmZl3d3d3d3d3d3dmZmZ3d3d3d3eIiIiZmZmZmZmqqqqqqqqqqqqqqqqqqqqqqqq7u7uqqqqqqqqqqqqZmZmZmZmIiIiIiIiIiIiIiIiIiIiZmZmIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3eIiIiIiIiqqqq7u7u7u7u7u7uqqqqZmZmIiIiIiIiIiIiZmZmZmZmIiIh3d3dmZmZmZmZmZmZ3d3eIiIiIiIiZmZmqqqqZmZmZmZmIiIiIiIh3d3d3d3eIiIiIiIiIiIiIiIiZmZmIiIiIiIh3d3d3d3dmZmZ3d3d3d3eIiIiZmZmqqqqZmZmIiIhmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3dmZmZVVVV3d3eIiIiqqqq7u7uqqqqqqqqZmZmZmZmZmZmZmZmIiIiIiIiIiIhmZmZVVVVVVVVmZmZmZmZmZmaIiIiZmZnMzMy7u7uqqqqZmZmIiIiIiIiqqqqqqqqqqqqZmZmZmZmqqqq7u7uqqqqZmZmqqqq7u7u7u7vMzMzMzMzMzMzMzMzMzMy7u7uqqqqZmZmIiIiIiIiIiIiIiIiIiIh3d3d3d3dmZmZ3d3eIiIiqqqqZmZl3d3d3d3eIiIiqqqq7u7u7u7vMzMy7u7u7u7uqqqqZmZmZmZmZmZmIiIiIiIh3d3d3d3dmZmZ3d3eIiIi7u7uqqqqqqqqIiIiIiIiIiIiqqqq7u7uZmZmIiIh3d3d3d3dmZmZmZmZ3d3eZmZmIiIiIiIh3d3eIiIiZmZmZmZmIiIh3d3dmZmZmZmaIiIiIiIh3d3d3d3dmZmZVVVVVVVVmZmaIiIh3d3eIiIiIiIiZmZmZmZmZmZmIiIhmZmZmZmZmZmZ3d3d3d3eqqqqZmZmZmZmIiIhVVVVmZmZmZmZ3d3dmZmZVVVVERERERERERERVVVVmZmZ3d3eIiIh3d3dmZmZmZmZmZmaIiIiIiIiIiIhmZmZmZmZmZmZmZmZmZmZ3d3d3d3eIiIiIiIiIiIiIiIiqqqq7u7u7u7uZmZmZmZmqqqq7u7vMzMzMzMy7u7u7u7uqqqrMzMy7u7uqqqqqqqq7u7u7u7u7u7uZmZmIiIiIiIi7u7uqqqqqqqq7u7uqqqqIiIiIiIiIiIiqqqqqqqqIiIiIiIiqqqq7u7vMzMzu7u7u7u7u7u7////u7u7////////u7u7MzMzMzMzd3d3///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3d3d3du7u7mZmZmZmZiIiImZmZqqqqmZmZmZmZiIiIiIiIiIiImZmZmZmZmZmZmZmZqqqqmZmZqqqqu7u7u7u7qqqqqqqqqqqqqqqqmZmZmZmZmZmZmZmZmZmZmZmZqqqqzMzM3d3dzMzMu7u7mZmZiIiId3d3ZmZmZmZmZmZmZmZmZmZmd3d3d3d3iIiId3d3iIiIiIiIiIiIiIiIiIiImZmZmZmZiIiIiIiId3d3d3d3ZmZmd3d3ZmZmd3d3iIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmd3d3iIiImZmZu7u7u7u7u7u7u7u7mZmZmZmZiIiIiIiIqqqqmZmZmZmZd3d3ZmZmVVVVVVVVd3d3d3d3iIiIiIiImZmZqqqqmZmZmZmZiIiId3d3iIiId3d3ZmZmd3d3d3d3d3d3iIiId3d3d3d3d3d3ZmZmd3d3d3d3mZmZqqqqqqqqmZmZiIiId3d3ZmZmZmZmd3d3d3d3d3d3d3d3ZmZmZmZmREREVVVVZmZmd3d3d3d3iIiImZmZmZmZmZmZmZmZmZmZmZmZmZmZd3d3ZmZmZmZmd3d3ZmZmZmZmZmZmd3d3mZmZu7u7zMzMqqqqmZmZiIiIiIiIqqqqu7u7qqqqmZmZmZmZu7u7u7u7qqqqmZmZqqqqqqqqu7u7u7u7zMzMzMzMzMzMzMzMzMzMu7u7qqqqiIiId3d3iIiImZmZmZmZiIiId3d3d3d3d3d3mZmZmZmZmZmZd3d3ZmZmiIiIqqqqzMzMzMzM3d3d3d3dzMzMzMzMqqqqmZmZiIiIiIiIiIiIiIiId3d3ZmZmd3d3mZmZu7u7qqqqqqqqiIiIiIiId3d3qqqqmZmZiIiIZmZmZmZmZmZmZmZmZmZmiIiIiIiIiIiId3d3ZmZmd3d3mZmZiIiIiIiId3d3ZmZmd3d3iIiId3d3d3d3ZmZmZmZmZmZmd3d3iIiImZmZiIiIiIiIiIiImZmZu7u7qqqqmQD//wAAmZl3d3dmZmZ3d3d3d3eIiIiZmZmqqqqZmZl3d3dmZmZVVVVmZmZ3d3dmZmZVVVVERERERERERERERERVVVVmZmZ3d3d3d3dmZmZmZmZ3d3eIiIiIiIh3d3d3d3dmZmZVVVVmZmZ3d3d3d3d3d3eIiIiIiIiqqqqZmZmZmZmqqqqqqqqZmZmZmZmqqqq7u7vMzMzMzMy7u7uqqqq7u7u7u7u7u7uqqqqqqqq7u7u7u7uqqqqIiIh3d3eIiIiqqqq7u7uqqqqqqqqqqqqIiIh3d3eIiIiqqqqqqqqIiIiIiIiqqqq7u7vd3d3d3d3u7u7u7u7u7u7u7u7MzMy7u7uZmZmqqqrMzMzu7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////7u7u////////////////////////////////////////////////7u7u7u7u3d3d7u7uzMzMqqqqmZmZmZmZqqqqqqqqmZmZiIiImZmZiIiIiIiIiIiImZmZmZmZqqqqqqqqmZmZqqqqqqqqqqqqqqqqu7u7u7u7qqqqu7u7qqqqmZmZiIiIiIiIiIiImZmZu7u7zMzM3d3d3d3du7u7qqqqiIiIZmZmZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmVVVVZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiImZmZu7u7zMzMu7u7u7u7mZmZiIiIiIiImZmZqqqqqqqqmZmZd3d3ZmZmVVVVVVVVZmZmd3d3iIiIiIiImZmZiIiImZmZmZmZmZmZiIiIiIiIZmZmd3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3ZmZmiIiImZmZqqqqqqqqmZmZiIiIZmZmZmZmZmZmd3d3d3d3iIiId3d3ZmZmVVVVREREREREVVVVVVVVZmZmd3d3d3d3mZmZmZmZmZmZiIiIiIiId3d3d3d3ZmZmd3d3ZmZmd3d3ZmZmd3d3iIiIqqqqu7u7u7u7qqqqqqqqmZmZqqqqqqqqu7u7qqqqiIiImZmZu7u7zMzMqqqqqqqqmZmZqqqqqqqqqqqqu7u7zMzMzMzMu7u7u7u7qqqqd3d3d3d3iIiIiIiImZmZiIiIiIiIiIiId3d3iIiIqqqqmZmZiIiId3d3iIiIqqqqzMzM3d3dzMzM3d3d3d3dzMzMzMzMqqqqmZmZmZmZiIiIiIiId3d3d3d3d3d3iIiIqqqqqqqqmZmZiIiId3d3d3d3iIiImZmZd3d3VVVVVVVVZmZmZmZmVVVVZmZmd3d3d3d3d3d3ZmZmd3d3iIiImZmZiIiIZmZmd3d3ZmZmZmZmZmZmd3d3ZmZmZmZmZmZmiIiIqqqqu7u7u7u7mZmZiIiImZmZqqqqqqqqqqqqiIiId3d3d3d3d3d3iIiIiIiIqqqqmZmZiIiIZmZmZmZmZmZmZmZmd3d3d3d3VVVVREREREREVVVVVVVVd3d3d3d3ZmZmZmZmZmZmd3d3d3d3mZmZiIiIZmZmVVVVVVVVZmZmZmZmd3d3d3d3d3d3mZmZmZmZqqqqqqqqqqqqqqqqmZmZmZmZmZmZu7u7zMzMzMzMqqqqqqqqu7u7u7u7u7u7qqqqqqqqmZmZu7u7qqqqiIiIZmZmZmZmmZmZqqqqqqqqiIiIiIiIiIiIZmZmd3d3mZmZu7u7qqqqqqqqqqqqu7u7zMzM3d3d7u7uzMzMu7u7zMzMzMzM3d3d3d3d3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7v///+7u7v///////////////////////+7u7t3d3czMzN3d3d3d3aqqqqqqqpmZmaqqqqqqqqqqqqqqqpmZmZmZmZmZmaqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqru7u7u7u6qqqqqqqqqqqqqqqqqqqqqqqpmZmYiIiIiIiIiIiJmZmaqqqszMzMzMzMzMzKqqqnd3d3d3d1VVVVVVVWZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZlVVVWZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiJmZmaqqqru7u8zMzLu7u6qqqpmZmYiIiIiIiJmZmYiIiIiIiIiIiFVVVVVVVVVVVVVVVXd3d2ZmZnd3d3d3d4iIiJmZmZmZmZmZmZmZmYiIiIiIiHd3d4iIiHd3d3d3d3d3d4iIiIiIiHd3d3d3d3d3d4iIiJmZmZmZmZmZmZmZmYiIiHd3d2ZmZnd3d3d3d4iIiIiIiHd3d2ZmZmZmZkRERFVVVVVVVVVVVVVVVWZmZnd3d4iIiIiIiIiIiIiIiJmZmYiIiGZmZnd3d3d3d3d3d3d3d2ZmZmZmZnd3d6qqqqqqqru7u7u7u6qqqpmZmZmZmbu7u7u7u6qqqoiIiKqqqru7u8zMzMzMzLu7u6qqqpmZmZmZmZmZmaqqqqqqqru7u7u7u6qqqpmZmYiIiHd3d4iIiJmZmZmZmZmZmYiIiHd3d3d3d4iIiJmZmZmZmXd3d3d3d4iIiLu7u93d3czMzN3d3d3d3d3d3d3d3czMzLu7u6qqqpmZmZmZmYiIiHd3d3d3d3d3d4iIiJmZmaqqqpmZmZmZmXd3d3d3d4iIiIiIiGZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZnd3d5mZmZmZmZmZmYiIiGZmZlVVVWZmZnd3d3d3d2ZmZmZmZnd3d5mZmaqqqru7u7u7u7u7u5mZmYiIiIiIiJmZmZmZmZmZmYiIiHd3d3d3d3d3d5mZmaqqqqqqqoiIiGZmZmZmZmZmZnd3d2ZmZmZmZlVVVURERERERFVVVWZmZnd3d3d3d3d3d3d3d2ZmZmZmZnd3d4iIiHd3d3d3d2ZmZmZmZmZmZnd3d3d3d3d3d3d3d5mZmbu7u6qqqqqqqqqqqru7u6qqqoiIiJmZmbu7u8zMzLu7u6qqqpmZmaqqqru7u6qqqqqqqpmZmYiIiJmZmaqqqpmZmXd3d3d3d4iIiIiIiHd3d3d3d3d3d2ZmZmZmZnd3d5mZmczMzLu7u7u7u6qqqru7u8zMzN3d3bu7u5mZmbu7u+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////u7u7////////u7u7////////////////u7u7////////////u7u7////////////////////////u7u7////////u7u7////////////////u7u7////////////////u7u7////////u7u7////////////u7u7////////u7u7d3d3d3d3u7u7u7u7u7u7////u7u7u7u7d3d3u7u7d3d3MzMzd3d3d3d3MzMzMzMzd3d3u7u7u7u7u7u7////////////d3d27u7vd3d3d3d27u7uqqqqZmZmZmZmqqqqqqqqqqqq7u7u7u7u7u7u7u7vMzMy7u7uqqqq7u7u7u7u7u7vMzMzMzMy7u7vMzMy7u7u7u7u7u7u7u7u7u7uqqqqqqqqqqqqIiIiIiIiIiIiqqqq7u7vMzMzMzMy7u7uZmZmIiIhmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZ3d3d3d3dmZmZmZmZ3d3dmZmZmZmZmZmZ3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmaIiIh3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiZmZm7u7u7u7u7u7u7u7uZmZmIiIh3d3d3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVVVVVmZmZmZmZ3d3d3d3eIiIiZmZmZmZmZmZmIiIiIiIiIiIiZmZmIiIiIiIh3d3eIiIiIiIiIiIh3d3d3d3d3d3eIiIiZmZmIiIiIiIiIiIiIiIiIiIhmZmZ3d3d3d3eIiIiIiIh3d3dmZmZVVVVVVVVERERVVVVVVVVVVVVmZmZ3d3d3d3d3d3eIiIiIiIh3d3dmZmZ3d3d3d3dmZmZmZmZmZmZ3d3d3d3eZmZm7u7u7u7u7u7uqqqqZmZmZmZm7u7vMzMyqqqqZmZmZmZm7u7vMzMzMzMzMzMy7u7uZmZmIiIiIiIiZmZmqqqq7u7u7u7uZmZmIiIh3d3d3d3eIiIiZmZmZmZmZmZmZmZmIiIiIiIiIiIiZmZmZmZmIiIh3d3eIiIi7u7vd3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMy7u7uqqqqZmZmIiIiIiIh3d3eIiIiIiIiZmZmqqqqqqqqIiIh3d3eIiIiIiIiIiIhmZmZmZmZ3d3eIiIh3d3d3d3dmZmZVVVVmZmZmZmZmZmZ3d3eZmZmZmZmqqqqIiIhmZmZVVVVVVVV3d3d3d3d3d3dmZmZmZmaIiIiqqqrMzMzMzMy7u7uZmZmIiIiIiIiZmZmZmZmIiIiIiIh3d3eIiIh3d3eZmZmZmZmqqqqIiIhmZmZmZmZmZmZmZmZmZmZVVVVVVVVERERVVVVmZmZmZmZ3d3eIiIiIiIh3d3dmZmZmZmZ3d3eIiIiIiIh3d3dmZmZmZmZmZmaIiIiIiIh3d3d3d3eZmZmqqqrMzMy7u7uqqqq7u7uqqqqIiIiIiIi7u7u7u7u7u7uZmZmIiIiZmZmqqqq7u7uZmZmIiIh3d3eZmZm7u7uqqqp3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZ3d3eZmZnMzMzMzMy7u7u7u7u7u7vMzMzMzMyqqqqqqqq7u7vd3d3////////////////////////////u7u7////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u3d3dzMzMu7u7mZmZiIiImZmZqqqqu7u7u7u73d3d3d3d3d3d3d3dzMzM3d3d3d3dzMzMzMzMqqqqqqqqu7u7u7u7zMzMzMzM3d3d7u7u3d3dzMzMu7u7zMzMqqqqqqqqqqqqqqqqqqqqu7u7qqqqu7u7u7u7zMzMzMzMzMzM3d3d3d3d3d3d7u7u3d3d3d3d3d3d3d3dzMzM3d3d3d3d3d3dzMzMzMzMu7u7zMzMu7u7qqqqmZmZiIiIiIiIiIiImZmZu7u7u7u7u7u7u7u7mZmZiIiId3d3ZmZmZmZmVVVVZmZmd3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmd3d3ZmZmd3d3ZmZmiIiId3d3d3d3iIiId3d3iIiIiIiId3d3iIiIiIiId3d3d3d3d3d3iIiIiIiImZmZu7u7u7u7u7u7qqqqiIiId3d3iIiId3d3d3d3iIiId3d3d3d3VVVVREREVVVVZmZmZmZmZmZmd3d3iIiImZmZiIiIiIiImZmZmZmZmZmZiIiImZmZiIiImZmZmZmZmZmZiIiIiIiIiIiId3d3d3d3iIiIiIiId3d3iIiId3d3ZmZmZmZmd3d3d3d3iIiIiIiIiIiIZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3iIiIiIiId3d3d3d3ZmZmVVVVZmZmZmZmZmZmd3d3mZmZqqqqzMzMqqqqqqqqqqqqmZmZu7u7zMzMu7u7mZmZiIiImZmZu7u7zMzMu7u7qqqqmZmZmZmZiIiIiIiImZmZmZmZmZmZmZmZiIiId3d3d3d3d3d3mZmZmZmZmZmZmZmZiIiIiIiIiIiImZmZqqqqiIiId3d3mZmZqqqq3d3d3d3dzMzM3d3d3d3d3d3dzMzM3d3du7u7qqqqmZmZiIiIiIiIiIiIiIiIiIiImZmZu7u7qqqqmZmZd3d3d3d3iIiIiIiId3d3ZmZmd3d3d3d3iIiId3d3ZmZmVVVVVVVVZmZmZmZmiIiIiIiIqqqqqqqqiIiIZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmiIiIqqqqu7u7u7u7u7u7qqqqmZmZiIiIiIiImZmZiIiIiIiIiIiId3d3iIiIiIiImZmZmZmZmZmZd3d3ZmZmd3d3iIiIiIiIZmZmREREVVVVZmZmiIiImZmZiIiIiIiImZmZiIiIZmZmZmZmd3d3iIiImZmZiIiId3d3ZmZmZmZmiIiIiIiId3d3d3d3iIiIqqqqzMzMu7u7u7u7qqqqmZmZiIiImZmZqqqqu7u7u7u7iIiIiIiIiIiImZmZmZmZiIiIZmZmd3d3qqqqu7u7u7u7iIiId3d3d3d3iIiId3d3d3d3ZmZmd3d3ZmZmZmZmiIiIzMzM3d3du7u7qqqqqqqqu7u7u7u7qqqqqqqqu7u7zMzM7u7u////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7t3d3d3d3d3d3bu7u6qqqqqqqoiIiHd3d3d3d4iIiIiIiJmZmZmZmZmZmaqqqqqqqszMzN3d3d3d3d3d3d3d3czMzMzMzKqqqqqqqqqqqqqqqqqqqqqqqru7u4iIiHd3d3d3d3d3d4iIiIiIiJmZmaqqqqqqqqqqqru7u7u7u8zMzO7u7u7u7u7u7u7u7v///+7u7v///+7u7u7u7u7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzLu7u6qqqpmZmYiIiHd3d4iIiKqqqqqqqru7u7u7u6qqqqqqqpmZmXd3d2ZmZlVVVWZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d4iIiIiIiJmZmZmZmZmZmZmZmZmZmYiIiJmZmZmZmZmZmZmZmYiIiIiIiIiIiIiIiHd3d4iIiIiIiKqqqqqqqru7u7u7u6qqqpmZmYiIiGZmZmZmZoiIiIiIiHd3d3d3d1VVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d5mZmYiIiJmZmaqqqpmZmaqqqqqqqqqqqqqqqpmZmZmZmYiIiIiIiHd3d3d3d4iIiIiIiHd3d3d3d2ZmZmZmZmZmZnd3d4iIiIiIiJmZmXd3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d4iIiJmZmXd3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d2ZmZoiIiKqqqqqqqru7u6qqqqqqqpmZmaqqqru7u8zMzJmZmXd3d3d3d6qqqqqqqqqqqqqqqqqqqpmZmXd3d4iIiHd3d4iIiHd3d3d3d3d3d3d3d2ZmZoiIiJmZmZmZmZmZmYiIiIiIiIiIiJmZmaqqqqqqqpmZmYiIiIiIiLu7u8zMzMzMzN3d3d3d3e7u7t3d3d3d3czMzMzMzLu7u6qqqoiIiJmZmYiIiHd3d4iIiJmZmaqqqru7u6qqqoiIiHd3d4iIiJmZmXd3d1VVVVVVVXd3d4iIiIiIiHd3d1VVVVVVVVVVVWZmZmZmZnd3d5mZmaqqqpmZmXd3d2ZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZoiIiKqqqqqqqszMzLu7u6qqqpmZmYiIiJmZmYiIiJmZmXd3d3d3d3d3d4iIiJmZmaqqqqqqqoiIiHd3d4iIiIiIiIiIiHd3d1VVVVVVVXd3d5mZmbu7u6qqqqqqqqqqqpmZmXd3d2ZmZnd3d4iIiJmZmYiIiGZmZmZmZmZmZnd3d3d3d3d3d2ZmZnd3d5mZmbu7u7u7u7u7u6qqqpmZmXd3d4iIiJmZmaqqqqqqqoiIiHd3d4iIiJmZmYiIiHd3d1VVVWZmZnd3d6qqqru7u5mZmXd3d3d3d4iIiIiIiGZmZmZmZmZmZmZmZmZmZnd3d7u7u93d3czMzKqqqpmZmaqqqqqqqqqqqqqqqpmZmZmZmd3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7d3d3d3d3d3d3MzMzMzMy7u7uqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqZmZmqqqqZmZm7u7u7u7vMzMzMzMzd3d3d3d3d3d3MzMzMzMzMzMyqqqqqqqqZmZmqqqp3d3dmZmZmZmZVVVVVVVVmZmZ3d3eIiIiIiIiqqqq7u7vMzMzMzMzd3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3MzMzMzMzMzMzMzMy7u7uqqqqqqqqZmZmIiIiIiIiIiIiZmZmZmZmqqqq7u7uqqqqIiIhmZmZmZmZmZmZVVVVmZmZVVVV3d3dmZmZmZmZmZmZVVVVmZmZ3d3eIiIiIiIiIiIiZmZmZmZmqqqqqqqqqqqqqqqq7u7uqqqq7u7uqqqqqqqq7u7uqqqqqqqqZmZmqqqqIiIiIiIh3d3eIiIiIiIiIiIiqqqq7u7u7u7u7u7uqqqqIiIh3d3dmZmZ3d3d3d3eIiIh3d3dmZmZVVVVERERVVVVVVVVmZmZVVVVmZmZ3d3d3d3eIiIiZmZmZmZmqqqq7u7uqqqq7u7u7u7u7u7u7u7uqqqqZmZmIiIiIiIh3d3eIiIiIiIiIiIiIiIiIiIh3d3dmZmaIiIiIiIiZmZmZmZmIiIhmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZ3d3dmZmZ3d3eIiIiZmZm7u7u7u7uZmZmZmZmIiIiZmZmqqqq7u7uIiIh3d3dmZmaIiIiZmZmZmZmZmZmZmZmIiIh3d3dmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3eZmZmZmZmZmZmIiIiIiIiZmZmZmZmqqqqZmZmZmZl3d3eIiIiqqqrMzMzMzMzd3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMyqqqqZmZmZmZmIiIh3d3eIiIiZmZm7u7uqqqqZmZl3d3d3d3eIiIiIiIhmZmZVVVVVVVVmZmZmZmZ3d3d3d3dmZmZVVVVVVVVmZmZmZmaIiIiqqqqqqqqIiIh3d3dmZmZmZmZ3d3d3d3d3d3d3d3dmZmZ3d3d3d3eZmZmZmZm7u7uqqqqqqqqqqqqZmZmZmZmIiIh3d3d3d3d3d3d3d3d3d3eqqqqqqqqqqqqZmZl3d3eIiIiIiIiZmZl3d3dmZmZmZmaIiIiZmZm7u7u7u7u7u7u7u7uqqqp3d3dmZmZ3d3eIiIiIiIh3d3dmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZ3d3eIiIiqqqq7u7u7u7uZmZmZmZl3d3d3d3eZmZmqqqqZmZl3d3d3d3d3d3eIiIiIiIhmZmZVVVVVVVV3d3eqqqqqqqqZmZl3d3dmZmZ3d3d3d3d3d3dmZmZ3d3dmZmZmZmZ3d3e7u7vMzMy7u7uqqqqZmZmqqqqqqqqqqqqZmZmIiIiIiIi7u7vu7u7////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////7u7u3d3dzMzM3d3d3d3d3d3du7u7u7u7u7u7u7u7u7u7zMzMzMzMzMzMzMzMu7u7zMzMu7u7u7u7u7u7qqqqu7u7qqqqqqqqzMzMzMzM3d3d3d3d3d3d3d3du7u7qqqqqqqqmZmZiIiIiIiId3d3ZmZmZmZmVVVVZmZmiIiImZmZqqqqu7u7u7u7u7u7u7u7zMzMzMzMzMzM3d3d3d3d7u7u3d3d3d3d7u7u3d3d3d3d3d3d3d3dzMzM3d3d3d3d3d3dzMzMzMzMu7u7zMzMu7u7qqqqiIiIiIiIiIiIiIiIiIiImZmZqqqqqqqqmZmZmZmZd3d3d3d3ZmZmZmZmVVVVVVVVZmZmd3d3d3d3ZmZmZmZmZmZmd3d3iIiIqqqqqqqqqqqqu7u7u7u7u7u7u7u7u7u7u7u7u7u7zMzMu7u7u7u7u7u7zMzMu7u7u7u7qqqqmZmZiIiIiIiIiIiIiIiId3d3iIiImZmZqqqqu7u7qqqqmZmZd3d3ZmZmZmZmd3d3d3d3d3d3d3d3ZmZmVVVVREREREREVVVVZmZmd3d3d3d3d3d3iIiImZmZqqqqu7u7u7u7u7u73d3dzMzM3d3du7u7u7u7qqqqmZmZiIiIiIiIiIiImZmZmZmZmZmZd3d3d3d3ZmZmiIiIiIiImZmZmZmZmZmZd3d3ZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmd3d3ZmZmd3d3iIiImZmZqqqqqqqqqqqqmZmZd3d3iIiImZmZmZmZiIiIZmZmZmZmZmZmd3d3d3d3mZmZiIiIiIiIZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3mZmZmZmZmZmZmZmZd3d3iIiIiIiImZmZmZmZiIiIiIiIiIiIqqqqzMzMzMzM7u7u3d3d3d3d3d3d3d3d3d3dzMzMzMzMu7u7mZmZmZmZiIiId3d3qqqqqqqqqqqqmZmZiIiId3d3d3d3iIiIiIiIZmZmVVVVREREREREVVVVd3d3d3d3ZmZmVVVVVVVVVVVVZmZmd3d3iIiIqqqqmZmZd3d3ZmZmZmZmZmZmiIiId3d3ZmZmVVVVd3d3d3d3iIiIiIiImZmZqqqqu7u7qqqqqqqqiIiIiIiId3d3d3d3ZmZmZmZmiIiIqqqqu7u7mZmZiIiId3d3iIiIqqqqqqqqmZmZd3d3d3d3mZmZqqqqu7u7u7u7zMzMzMzMu7u7mZmZd3d3ZmZmiIiIiIiId3d3ZmZmZmZmd3d3d3d3d3d3ZmZmZmZmd3d3mZmZqqqqu7u7qqqqiIiId3d3d3d3iIiIiIiImZmZqqqqiIiId3d3iIiImZmZiIiIZmZmVVVVVVVVZmZmmZmZu7u7mZmZiIiIZmZmiIiId3d3ZmZmd3d3d3d3ZmZmVVVVd3d3mZmZu7u7zMzMqqqqmZmZqqqqu7u7qqqqiIiId3d3iIiIqqqq3d3d////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////+7u7v///////////////////////////////////////////////////////+7u7v///////////////////+7u7t3d3czMzLu7u8zMzMzMzN3d3czMzMzMzMzMzN3d3d3d3d3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3czMzLu7u6qqqoiIiIiIiIiIiKqqqszMzN3d3d3d3d3d3czMzLu7u7u7u6qqqqqqqqqqqpmZmYiIiHd3d3d3d3d3d3d3d4iIiJmZmZmZmaqqqru7u8zMzMzMzMzMzN3d3d3d3d3d3e7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7t3d3d3d3czMzLu7u8zMzLu7u6qqqpmZmYiIiHd3d3d3d4iIiIiIiJmZmaqqqqqqqqqqqoiIiHd3d3d3d2ZmZmZmZlVVVWZmZnd3d3d3d3d3d3d3d3d3d3d3d4iIiKqqqqqqqru7u7u7u6qqqru7u8zMzMzMzLu7u8zMzMzMzLu7u8zMzMzMzLu7u8zMzLu7u6qqqqqqqqqqqpmZmYiIiIiIiHd3d4iIiJmZmZmZmbu7u7u7u6qqqoiIiHd3d2ZmZmZmZnd3d3d3d3d3d3d3d2ZmZlVVVVVVVWZmZoiIiIiIiIiIiIiIiJmZmaqqqqqqqru7u8zMzMzMzN3d3d3d3czMzMzMzLu7u7u7u6qqqpmZmZmZmZmZmZmZmZmZmZmZmXd3d3d3d3d3d3d3d3d3d4iIiKqqqpmZmXd3d2ZmZlVVVVVVVWZmZmZmZlVVVVVVVWZmZmZmZnd3d2ZmZnd3d2ZmZnd3d2ZmZnd3d3d3d3d3d4iIiHd3d3d3d4iIiKqqqqqqqpmZmYiIiHd3d3d3d4iIiJmZmZmZmXd3d0RERFVVVVVVVWZmZnd3d4iIiGZmZmZmZnd3d2ZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZoiIiJmZmZmZmYiIiIiIiHd3d4iIiIiIiJmZmZmZmXd3d3d3d5mZmbu7u8zMzMzMzMzMzN3d3d3d3czMzN3d3d3d3czMzLu7u5mZmYiIiIiIiKqqqqqqqpmZmZmZmZmZmYiIiHd3d3d3d3d3d3d3d3d3d1VVVURERERERFVVVXd3d3d3d3d3d2ZmZlVVVVVVVWZmZnd3d5mZmaqqqpmZmXd3d2ZmZmZmZnd3d4iIiIiIiGZmZmZmZnd3d4iIiJmZmZmZmYiIiKqqqru7u7u7u6qqqqqqqoiIiIiIiIiIiHd3d3d3d4iIiJmZmZmZmZmZmYiIiHd3d4iIiKqqqru7u5mZmXd3d4iIiJmZmbu7u7u7u7u7u7u7u8zMzMzMzJmZmXd3d3d3d5mZmYiIiHd3d3d3d2ZmZmZmZoiIiHd3d3d3d2ZmZmZmZoiIiKqqqqqqqqqqqpmZmXd3d3d3d3d3d4iIiKqqqqqqqoiIiHd3d4iIiJmZmZmZmXd3d2ZmZlVVVWZmZqqqqru7u5mZmYiIiHd3d4iIiIiIiGZmZnd3d4iIiGZmZmZmZmZmZoiIiKqqqszMzKqqqpmZmaqqqru7u6qqqqqqqoiIiHd3d5mZmd3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7u7u7u7u7////////////////u7u7////////////////////////////////////////////////////u7u7////////////////u7u7u7u7u7u7u7u7u7u7u7u7////////////////////////d3d27u7u7u7uqqqqqqqrMzMzMzMzd3d3MzMzd3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3MzMy7u7uIiIiIiIiIiIiIiIiIiIiZmZmqqqrMzMzMzMy7u7u7u7u7u7u7u7uqqqq7u7uqqqqZmZmIiIh3d3d3d3d3d3d3d3eIiIiIiIiZmZmqqqq7u7vMzMzMzMzd3d3d3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3u7u7d3d3MzMzMzMy7u7u7u7u7u7uqqqqqqqqIiIiIiIh3d3d3d3eIiIiZmZmZmZmZmZmZmZmZmZmZmZmIiIh3d3d3d3dmZmZmZmZ3d3d3d3d3d3d3d3eIiIh3d3eIiIiZmZmqqqq7u7u7u7vMzMy7u7vMzMy7u7u7u7u7u7vMzMy7u7vMzMy7u7vMzMy7u7u7u7uqqqqqqqqqqqqZmZmIiIh3d3eIiIh3d3eIiIiZmZmZmZmqqqqqqqqZmZl3d3d3d3dmZmZmZmZ3d3eIiIiIiIh3d3dmZmZmZmZ3d3d3d3eZmZmqqqq7u7uqqqqqqqq7u7u7u7u7u7vMzMzMzMzMzMzMzMzMzMy7u7u7u7uqqqqZmZmIiIiIiIiIiIiZmZmZmZmIiIiIiIhmZmZmZmZ3d3eZmZmZmZmqqqqIiIhmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3dmZmZ3d3d3d3eIiIiIiIiIiIiIiIiIiIh3d3eIiIiIiIiqqqqZmZmZmZmIiIh3d3eIiIiqqqqZmZl3d3dERERVVVVVVVVmZmZ3d3d3d3d3d3d3d3eIiIh3d3dmZmZVVVVmZmZVVVVmZmZmZmZmZmaIiIiqqqqZmZmZmZmIiIh3d3d3d3eIiIiqqqqZmZl3d3dmZmaZmZm7u7vMzMzMzMzMzMzMzMzd3d3d3d3d3d3d3d3MzMy7u7uZmZmIiIiIiIiIiIh3d3d3d3eZmZmZmZmZmZl3d3d3d3d3d3eIiIhmZmZVVVVERERVVVVVVVVmZmZ3d3d3d3d3d3dmZmZmZmZ3d3d3d3eZmZmZmZmZmZmIiIhmZmZmZmZ3d3eIiIiZmZl3d3d3d3eIiIiZmZmqqqqZmZmIiIiZmZmZmZm7u7u7u7u7u7uZmZmIiIiIiIh3d3d3d3d3d3eZmZmZmZmqqqqZmZmIiIiIiIiqqqq7u7uqqqp3d3eIiIiqqqq7u7u7u7u7u7uqqqq7u7u7u7uZmZl3d3eIiIiZmZmIiIiIiIhmZmZ3d3eIiIiIiIiIiIh3d3dmZmZ3d3eIiIiqqqqqqqqqqqqZmZl3d3dmZmZ3d3eIiIiqqqqqqqqIiIh3d3eIiIiZmZmZmZlmZmZmZmZVVVV3d3eqqqq7u7uqqqp3d3d3d3eIiIiIiIh3d3d3d3d3d3dmZmZmZmZmZmZ3d3eqqqq7u7uqqqqIiIiZmZm7u7u7u7uqqqqIiIh3d3eIiIjMzMzu7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u3d3d3d3d3d3d3d3d3d3d7u7u7u7u////7u7u////7u7u////////7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d7u7u////7u7u7u7u7u7uzMzMzMzMzMzM3d3d3d3d3d3d7u7u7u7u7u7u////u7u7iIiImZmZqqqqzMzMzMzMzMzMu7u7u7u7u7u7zMzMzMzM7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3dzMzMmZmZmZmZiIiIiIiImZmZiIiId3d3mZmZmZmZqqqqqqqqu7u7u7u7u7u7u7u7zMzMu7u7qqqqqqqqiIiIiIiIiIiIiIiImZmZiIiImZmZmZmZmZmZu7u7zMzMzMzM3d3dzMzM3d3d3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d3d3du7u7u7u7u7u7mZmZqqqqqqqqmZmZiIiIiIiId3d3d3d3iIiId3d3iIiImZmZmZmZqqqqmZmZmZmZmZmZd3d3d3d3ZmZmZmZmZmZmd3d3iIiIiIiIiIiIiIiImZmZqqqqu7u7qqqqzMzMu7u7u7u7u7u7u7u7zMzMzMzMu7u7zMzMu7u7zMzMu7u7u7u7u7u7u7u7qqqqmZmZiIiId3d3d3d3iIiIiIiId3d3iIiIqqqqu7u7u7u7mZmZd3d3d3d3ZmZmd3d3d3d3iIiImZmZd3d3ZmZmd3d3mZmZu7u7u7u7zMzMu7u7u7u7u7u7u7u7u7u7zMzMzMzMzMzMzMzMu7u7u7u7u7u7qqqqmZmZiIiId3d3iIiImZmZmZmZiIiId3d3d3d3ZmZmd3d3iIiImZmZqqqqiIiIZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3iIiImZmZiIiIiIiIiIiImZmZmZmZiIiImZmZqqqqqqqqmZmZiIiId3d3iIiIqqqqiIiIZmZmVVVVREREZmZmd3d3d3d3d3d3iIiIiIiId3d3d3d3ZmZmVVVVVVVVZmZmZmZmZmZmd3d3iIiIqqqqmZmZiIiIiIiId3d3iIiImZmZmZmZiIiId3d3d3d3mZmZqqqqzMzMzMzM3d3d3d3d3d3d3d3d3d3dzMzMzMzMqqqqmZmZd3d3d3d3ZmZmd3d3mZmZqqqqqqqqiIiIiIiId3d3d3d3iIiIZmZmVVVVVVVVZmZmd3d3d3d3iIiIiIiId3d3ZmZmZmZmZmZmd3d3mZmZqqqqqqqqiIiId3d3ZmZmiIiImZmZiIiId3d3ZmZmiIiIqqqqqqqqqqqqmZmZmZmZqqqqqqqqu7u7qqqqmZmZiIiId3d3d3d3ZmZmd3d3mZmZu7u7qqqqmZmZd3d3iIiIu7u7u7u7qqqqiIiId3d3qqqqu7u7zMzMu7u7qqqqqqqqqqqqmZmZiIiId3d3mZmZiIiIiIiId3d3d3d3qqqqmZmZmZmZd3d3ZmZmd3d3mZmZqqqqqqqqqqqqqqqqd3d3d3d3ZmZmiIiIu7u7mZmZiIiId3d3iIiImZmZiIiIZmZmVVVVZmZmiIiIu7u7u7u7qqqqiIiIiIiId3d3d3d3iIiId3d3iIiId3d3ZmZmZmZmd3d3iIiImZmZmZmZiIiImZmZqqqqu7u7qqqqiIiId3d3iIiIqqqq7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////+7u7v///////////+7u7v///////////////////+7u7v///////////////+7u7v///////+7u7v///////////////////////////////////////////+7u7v///////+7u7v///+7u7u7u7u7u7u7u7v///+7u7v///////////////+7u7t3d3d3d3czMzMzMzN3d3e7u7t3d3d3d3d3d3d3d3czMzMzMzN3d3czMzN3d3d3d3d3d3czMzMzMzLu7u7u7u7u7u8zMzN3d3d3d3e7u7u7u7t3d3d3d3czMzMzMzLu7u6qqqqqqqru7u8zMzMzMzJmZmWZmZmZmZqqqqru7u7u7u7u7u5mZmYiIiKqqqqqqqszMzN3d3d3d3d3d3e7u7u7u7u7u7u7u7u7u7szMzKqqqpmZmZmZmZmZmYiIiIiIiHd3d3d3d3d3d3d3d2ZmZnd3d4iIiJmZmaqqqru7u8zMzMzMzMzMzLu7u7u7u6qqqpmZmaqqqqqqqpmZmZmZmZmZmZmZmZmZmZmZmaqqqqqqqru7u8zMzMzMzMzMzN3d3d3d3d3d3d3d3d3d3czMzN3d3czMzMzMzMzMzLu7u7u7u6qqqpmZmZmZmZmZmZmZmZmZmYiIiIiIiHd3d3d3d4iIiIiIiHd3d4iIiJmZmaqqqqqqqqqqqpmZmYiIiHd3d3d3d2ZmZmZmZmZmZoiIiIiIiIiIiIiIiIiIiJmZmZmZmbu7u7u7u7u7u7u7u8zMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u6qqqpmZmYiIiHd3d3d3d3d3d4iIiHd3d4iIiJmZmaqqqru7u5mZmZmZmXd3d2ZmZmZmZnd3d5mZmaqqqpmZmYiIiIiIiJmZmbu7u7u7u8zMzMzMzLu7u7u7u7u7u7u7u7u7u8zMzLu7u8zMzLu7u7u7u7u7u7u7u5mZmZmZmYiIiIiIiIiIiIiIiJmZmYiIiGZmZlVVVWZmZoiIiJmZmaqqqpmZmXd3d1VVVVVVVVVVVWZmZmZmZnd3d2ZmZmZmZnd3d3d3d3d3d3d3d4iIiIiIiJmZmZmZmZmZmaqqqqqqqpmZmZmZmZmZmaqqqqqqqpmZmXd3d3d3d4iIiIiIiHd3d3d3d0RERERERFVVVWZmZnd3d4iIiHd3d3d3d3d3d2ZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZoiIiJmZmZmZmZmZmYiIiHd3d4iIiKqqqqqqqpmZmYiIiHd3d4iIiKqqqt3d3czMzN3d3d3d3czMzN3d3d3d3bu7u7u7u6qqqoiIiHd3d2ZmZnd3d4iIiIiIiJmZmZmZmYiIiHd3d3d3d4iIiIiIiIiIiFVVVVVVVXd3d3d3d3d3d5mZmZmZmZmZmXd3d3d3d2ZmZnd3d4iIiJmZmZmZmZmZmXd3d2ZmZnd3d4iIiJmZmXd3d3d3d3d3d5mZmbu7u7u7u7u7u7u7u6qqqqqqqqqqqqqqqqqqqoiIiHd3d2ZmZmZmZoiIiJmZmaqqqqqqqoiIiIiIiJmZmbu7u7u7u6qqqnd3d4iIiJmZmczMzMzMzMzMzKqqqqqqqqqqqpmZmYiIiHd3d5mZmZmZmYiIiIiIiIiIiJmZmZmZmZmZmXd3d3d3d3d3d6qqqqqqqqqqqqqqqqqqqnd3d2ZmZmZmZoiIiKqqqru7u4iIiGZmZnd3d5mZmZmZmXd3d1VVVVVVVXd3d5mZmaqqqpmZmXd3d3d3d3d3d4iIiIiIiIiIiHd3d2ZmZmZmZmZmZmZmZmZmZoiIiHd3d3d3d4iIiJmZmaqqqqqqqoiIiGZmZnd3d5mZmd3d3e7u7v///////+7u7v///////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////u7u7////////////u7u7////u7u7d3d3u7u7d3d3d3d3MzMy7u7uqqqqZmZmqqqq7u7vMzMzd3d3d3d3u7u7////////////u7u7u7u7u7u7d3d3u7u7d3d3MzMy7u7uqqqqqqqqZmZmZmZmqqqqqqqq7u7u7u7vMzMy7u7u7u7u7u7u7u7uZmZmqqqqZmZmqqqq7u7vMzMzMzMzd3d3d3d3d3d27u7uqqqqZmZmqqqqZmZmZmZl3d3eIiIiIiIh3d3eIiIiZmZmZmZmZmZmIiIiqqqq7u7u7u7vd3d3d3d3d3d3d3d3u7u7d3d3d3d3MzMyqqqqqqqqqqqqqqqqqqqqZmZmIiIiIiIiIiIh3d3dmZmZmZmZVVVVmZmaIiIiZmZmqqqrMzMzMzMzd3d3MzMzMzMzMzMy7u7uqqqqqqqqZmZmZmZmqqqqqqqqqqqqZmZmZmZmqqqqqqqqqqqq7u7vMzMy7u7vMzMzMzMzMzMzMzMzMzMy7u7vMzMy7u7uqqqqqqqqqqqqZmZmIiIiZmZmIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIiIiIiZmZmqqqqqqqqqqqqZmZmIiIh3d3d3d3dmZmZ3d3d3d3eIiIiIiIiIiIiZmZmIiIiZmZmqqqqqqqq7u7u7u7u7u7vd3d3MzMzMzMzMzMzMzMzd3d3MzMy7u7uqqqqqqqqqqqqqqqqZmZmZmZmIiIh3d3d3d3d3d3d3d3d3d3eIiIiZmZm7u7uqqqqqqqqZmZmIiIh3d3d3d3eZmZmqqqqqqqqZmZmIiIiIiIiqqqqqqqq7u7vMzMzd3d3d3d3MzMy7u7u7u7u7u7u7u7vMzMy7u7uqqqq7u7u7u7u7u7uZmZlmZmZ3d3d3d3eIiIiIiIh3d3d3d3dmZmZmZmZmZmaZmZmqqqqqqqqIiIhmZmZVVVVVVVVmZmZmZmZ3d3dmZmZ3d3eIiIiIiIh3d3eIiIiIiIiZmZmZmZmZmZmqqqqqqqq7u7uqqqqZmZmqqqqZmZmZmZmIiIiIiIh3d3dmZmZ3d3eIiIhmZmZERERERERVVVVmZmZ3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZ3d3eIiIiZmZmIiIh3d3eIiIiIiIiqqqqqqqqZmZmIiIh3d3eIiIiqqqrMzMzMzMzMzMzd3d3MzMzMzMy7u7uqqqqqqqqZmZl3d3d3d3d3d3d3d3d3d3eIiIiZmZmZmZl3d3dmZmZ3d3eIiIiZmZmIiIh3d3d3d3eIiIiZmZmIiIiZmZmqqqqqqqqIiIh3d3dmZmZ3d3d3d3eIiIiZmZmIiIh3d3dmZmZ3d3eIiIiZmZl3d3dmZmZ3d3eqqqq7u7vd3d3d3d3MzMy7u7uqqqqqqqqZmZmZmZmIiIh3d3dmZmZ3d3d3d3eZmZmqqqqqqqqZmZl3d3eIiIi7u7u7u7uZmZmIiIh3d3eZmZm7u7vMzMzMzMy7u7uqqqqqqqqIiIiIiIiIiIiZmZmZmZmIiIh3d3d3d3eIiIiZmZmIiIh3d3d3d3eIiIi7u7uqqqqqqqqZmZmZmZl3d3d3d3dmZmaIiIiqqqq7u7uIiIh3d3dmZmaZmZmIiIh3d3dVVVVVVVVVVVWIiIiZmZmZmZl3d3dmZmZ3d3eZmZmIiIh3d3dmZmZVVVVmZmZmZmZVVVVmZmZmZmZmZmZmZmZ3d3eZmZmqqqqZmZmZmZlmZmZmZmZ3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u3d3dzMzMu7u7zMzMzMzMu7u7qqqqmZmZiIiIiIiId3d3iIiImZmZqqqqu7u7zMzM3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7uzMzMzMzMu7u7u7u7qqqqiIiIiIiIiIiIiIiImZmZmZmZqqqqqqqqqqqqqqqqmZmZiIiIiIiId3d3iIiIiIiImZmZu7u7u7u7zMzMzMzMu7u7u7u7u7u7qqqqqqqqqqqqmZmZiIiIiIiIiIiIiIiImZmZiIiIiIiIiIiIiIiImZmZmZmZqqqqu7u7zMzMzMzM3d3dzMzMzMzMu7u7u7u7zMzMqqqqqqqqmZmZmZmZmZmZmZmZiIiImZmZd3d3ZmZmZmZmZmZmd3d3iIiImZmZqqqqzMzMzMzMzMzM3d3dzMzMu7u7u7u7qqqqqqqqmZmZqqqqu7u7u7u7qqqqqqqqqqqqmZmZqqqqmZmZmZmZqqqqzMzMzMzMu7u7u7u7u7u7zMzMu7u7u7u7qqqqmZmZmZmZmZmZiIiIiIiIiIiIiIiId3d3mZmZmZmZmZmZiIiId3d3iIiId3d3iIiId3d3iIiImZmZqqqqqqqqmZmZiIiId3d3d3d3iIiId3d3d3d3d3d3iIiIiIiImZmZmZmZmZmZmZmZqqqqqqqqu7u7u7u7zMzMu7u7zMzMzMzMu7u7zMzMzMzMu7u7u7u7qqqqmZmZmZmZiIiIiIiId3d3d3d3d3d3ZmZmd3d3ZmZmd3d3iIiImZmZu7u7qqqqmZmZiIiId3d3iIiIiIiIqqqqqqqqqqqqmZmZmZmZiIiIqqqqzMzM3d3dzMzM3d3dzMzMzMzMzMzMu7u7u7u7u7u7qqqqu7u7u7u7u7u7qqqqiIiId3d3ZmZmd3d3iIiIiIiId3d3ZmZmZmZmZmZmZmZmiIiImZmZmZmZiIiIZmZmREREVVVVZmZmd3d3d3d3iIiImZmZmZmZiIiImZmZmZmZmZmZiIiIqqqqqqqqqqqqu7u7qqqqqqqqmZmZmZmZmZmZmZmZmZmZmZmZd3d3ZmZmd3d3iIiIZmZmVVVVVVVVVVVVZmZmZmZmZmZmd3d3iIiId3d3d3d3d3d3ZmZmZmZmd3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiId3d3iIiIiIiIqqqqmZmZiIiIZmZmd3d3mZmZu7u7zMzMzMzMzMzMzMzMu7u7qqqqmZmZmZmZiIiId3d3d3d3ZmZmZmZmd3d3mZmZmZmZiIiIiIiId3d3ZmZmiIiImZmZiIiIZmZmd3d3mZmZmZmZmZmZqqqqu7u7qqqqmZmZiIiId3d3d3d3ZmZmiIiImZmZd3d3d3d3ZmZmd3d3iIiImZmZiIiIZmZmd3d3qqqqu7u7zMzMzMzMzMzMu7u7qqqqmZmZiIiId3d3ZmZmZmZmZmZmZmZmiIiImZmZqqqqqqqqiIiIiIiIiIiIqqqqu7u7mZmZd3d3d3d3iIiIqqqqu7u7zMzMu7u7u7u7qqqqiIiId3d3iIiIiIiIiIiIiIiId3d3d3d3iIiIiIiIiIiId3d3d3d3iIiIu7u7qqqqmZmZiIiIiIiId3d3ZmZmd3d3mZmZqqqqqqqqiIiIZmZmd3d3iIiIiIiId3d3VVVVREREZmZmZmZmd3d3d3d3ZmZmZmZmd3d3d3d3ZmZmZmZmVVVVVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVZmZmiIiImZmZqqqqiIiId3d3ZmZmd3d3u7u77u7u////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////+7u7t3d3d3d3e7u7t3d3czMzMzMzLu7u7u7u7u7u6qqqru7u6qqqpmZmZmZmYiIiIiIiJmZmZmZmZmZmZmZmbu7u7u7u8zMzMzMzN3d3e7u7u7u7t3d3czMzMzMzN3d3d3d3czMzMzMzKqqqqqqqoiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d6qqqru7u7u7u8zMzMzMzMzMzMzMzLu7u7u7u6qqqpmZmYiIiIiIiJmZmYiIiIiIiHd3d2ZmZmZmZnd3d2ZmZoiIiJmZmbu7u7u7u8zMzMzMzLu7u6qqqqqqqpmZmaqqqqqqqpmZmZmZmZmZmZmZmYiIiIiIiIiIiIiIiIiIiHd3d3d3d4iIiIiIiJmZmbu7u7u7u8zMzN3d3czMzMzMzLu7u7u7u7u7u6qqqqqqqqqqqru7u7u7u6qqqru7u6qqqoiIiIiIiIiIiKqqqru7u6qqqqqqqqqqqqqqqqqqqqqqqpmZmZmZmZmZmYiIiIiIiIiIiHd3d3d3d3d3d4iIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d2ZmZnd3d3d3d3d3d5mZmZmZmZmZmZmZmYiIiIiIiHd3d3d3d3d3d3d3d3d3d4iIiJmZmZmZmZmZmZmZmaqqqqqqqru7u6qqqru7u8zMzMzMzLu7u8zMzLu7u7u7u7u7u7u7u6qqqpmZmYiIiIiIiGZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZnd3d5mZmbu7u7u7u6qqqpmZmZmZmZmZmYiIiJmZmaqqqru7u6qqqpmZmZmZmZmZmbu7u7u7u8zMzN3d3d3d3czMzN3d3czMzLu7u7u7u6qqqru7u6qqqqqqqpmZmYiIiHd3d2ZmZmZmZmZmZoiIiHd3d3d3d3d3d2ZmZmZmZnd3d6qqqqqqqqqqqoiIiFVVVVVVVWZmZoiIiIiIiJmZmaqqqqqqqpmZmaqqqpmZmZmZmZmZmaqqqqqqqqqqqru7u6qqqpmZmZmZmZmZmaqqqru7u6qqqnd3d2ZmZlVVVWZmZnd3d2ZmZmZmZkRERFVVVVVVVVVVVWZmZmZmZnd3d3d3d4iIiHd3d3d3d4iIiHd3d4iIiGZmZnd3d3d3d4iIiJmZmXd3d2ZmZnd3d2ZmZpmZmaqqqoiIiHd3d2ZmZmZmZnd3d6qqqqqqqru7u7u7u6qqqqqqqqqqqoiIiJmZmYiIiHd3d3d3d2ZmZnd3d3d3d3d3d5mZmYiIiHd3d2ZmZmZmZnd3d4iIiIiIiGZmZnd3d6qqqqqqqqqqqpmZmbu7u8zMzKqqqpmZmXd3d3d3d3d3d4iIiIiIiIiIiHd3d2ZmZnd3d3d3d4iIiIiIiGZmZnd3d4iIiJmZmaqqqru7u7u7u6qqqpmZmYiIiHd3d2ZmZlVVVVVVVVVVVXd3d5mZmZmZmaqqqoiIiIiIiHd3d4iIiJmZmbu7u5mZmXd3d3d3d4iIiJmZmaqqqru7u8zMzLu7u6qqqoiIiHd3d3d3d4iIiIiIiIiIiGZmZnd3d3d3d4iIiHd3d2ZmZnd3d4iIiKqqqqqqqqqqqoiIiHd3d3d3d2ZmZnd3d5mZmaqqqpmZmXd3d2ZmZnd3d4iIiJmZmXd3d1VVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZnd3d4iIiJmZmZmZmXd3d2ZmZoiIiMzMzP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////u7u7u7u7u7u7u7u7u7u7d3d3MzMy7u7u7u7u7u7uqqqq7u7u7u7uqqqqqqqqqqqqIiIiZmZmZmZmZmZmIiIiIiIiIiIiIiIiZmZmZmZmqqqqqqqqqqqrMzMzd3d3u7u7u7u7u7u7u7u7d3d3MzMyqqqqqqqqqqqqZmZmZmZmIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmaIiIiZmZmZmZm7u7vMzMzMzMzMzMzMzMzMzMy7u7uqqqqqqqqqqqqZmZmIiIh3d3dmZmZ3d3d3d3d3d3d3d3eIiIiIiIiqqqq7u7u7u7uZmZl3d3d3d3eIiIiIiIiIiIiZmZmIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIiIiIiIiIiIiIiIiIiZmZmZmZm7u7u7u7vMzMzMzMzMzMzd3d3MzMy7u7uqqqqqqqqqqqqqqqq7u7u7u7u7u7uqqqqqqqqqqqqZmZmIiIiIiIh3d3d3d3d3d3eIiIiIiIiIiIiZmZl3d3eIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3eIiIiZmZmqqqqZmZmIiIiIiIiIiIh3d3dmZmZ3d3d3d3eIiIiZmZmqqqqqqqqZmZmZmZmZmZmZmZmqqqqqqqqqqqq7u7uqqqqqqqqqqqqZmZmqqqqqqqqZmZmZmZmIiIhmZmZVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmZ3d3eZmZmqqqq7u7u7u7uqqqqqqqqZmZmZmZmqqqq7u7u7u7uqqqqZmZmIiIiZmZmqqqrMzMzMzMzd3d3d3d3d3d3MzMy7u7uqqqqqqqqqqqqZmZmZmZmZmZmIiIh3d3dmZmZmZmZmZmZ3d3eIiIh3d3d3d3dmZmZmZmZ3d3eZmZmqqqqqqqqIiIhVVVVmZmaIiIiIiIiZmZmqqqqqqqqqqqqZmZmZmZmZmZmqqqqqqqqqqqqqqqqqqqqqqqq7u7uqqqqZmZmZmZmqqqqqqqqIiIiIiIhmZmZVVVVmZmZmZmZmZmZVVVVERERERERmZmZmZmZmZmZ3d3eIiIiZmZmZmZl3d3d3d3d3d3d3d3eIiIh3d3dmZmZ3d3d3d3eIiIiIiIh3d3dmZmZ3d3eZmZmZmZmZmZl3d3dmZmZVVVVmZmZ3d3eIiIiZmZmZmZmqqqqqqqqZmZmIiIiIiIh3d3d3d3dmZmZmZmZ3d3d3d3eIiIiZmZmIiIh3d3dmZmZmZmZmZmZ3d3dmZmZmZmZ3d3eZmZmqqqq7u7u7u7vMzMzMzMzMzMyZmZmIiIhmZmZ3d3eIiIiIiIiIiIhmZmZmZmZmZmZ3d3eIiIh3d3dmZmZmZmZmZmZ3d3eZmZmZmZmZmZmIiIiIiIiIiIh3d3dmZmZmZmZVVVVmZmZ3d3eIiIiqqqqZmZmIiIh3d3d3d3eIiIiZmZm7u7uZmZl3d3dmZmZ3d3eZmZm7u7u7u7u7u7u7u7u7u7uZmZl3d3d3d3d3d3eIiIhmZmZmZmZ3d3eIiIh3d3d3d3d3d3dmZmZ3d3e7u7uqqqqZmZmIiIh3d3dmZmZmZmZ3d3eZmZmZmZmZmZl3d3dmZmaIiIiZmZmIiIhmZmZVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZmZmZ3d3d3d3dmZmZmZmZmZmZ3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVV3d3eIiIiqqqqqqqqIiIhmZmaIiIjMzMzu7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////7u7u////7u7u////////////////////////7u7u7u7u7u7u7u7u////7u7u////7u7u7u7u7u7u7u7u7u7u////7u7u3d3dzMzM3d3d3d3d3d3d3d3dzMzMu7u7u7u7zMzMu7u7zMzMu7u7u7u7qqqqu7u7qqqqu7u7qqqqqqqqqqqqmZmZiIiId3d3d3d3iIiIiIiIiIiImZmZmZmZqqqqzMzM3d3d7u7u7u7u7u7u3d3dzMzMzMzMu7u7mZmZiIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3iIiIiIiImZmZu7u7zMzMzMzMzMzM3d3dzMzMu7u7u7u7u7u7mZmZiIiIiIiImZmZiIiIiIiImZmZiIiIiIiIiIiIiIiIiIiIZmZmREREREREVVVVZmZmZmZmd3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiId3d3iIiIiIiIiIiImZmZiIiImZmZmZmZu7u7zMzMzMzM3d3dzMzM3d3du7u7u7u7qqqqu7u7qqqqu7u7zMzMzMzMzMzMqqqqqqqqd3d3d3d3d3d3ZmZmZmZmZmZmd3d3ZmZmd3d3d3d3iIiIiIiIiIiId3d3iIiId3d3d3d3d3d3iIiId3d3iIiId3d3d3d3d3d3d3d3ZmZmZmZmZmZmiIiIiIiImZmZmZmZmZmZmZmZiIiId3d3d3d3d3d3d3d3iIiImZmZmZmZqqqqmZmZmZmZiIiIiIiIiIiIiIiImZmZiIiIiIiId3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiId3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3iIiIqqqqu7u7u7u7u7u7qqqqqqqqmZmZu7u7u7u7u7u7u7u7qqqqmZmZmZmZqqqqu7u7zMzMzMzMzMzMzMzMu7u7qqqqqqqqqqqqmZmZmZmZmZmZiIiId3d3d3d3ZmZmZmZmd3d3d3d3d3d3d3d3ZmZmZmZmVVVVd3d3iIiIqqqqqqqqiIiIZmZmZmZmiIiImZmZqqqqqqqqu7u7qqqqqqqqqqqqqqqqqqqqqqqqu7u7qqqqqqqqqqqqu7u7qqqqmZmZqqqqmZmZmZmZiIiId3d3ZmZmVVVVVVVVZmZmVVVVVVVVVVVVVVVVZmZmd3d3iIiIiIiIqqqqqqqqd3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3iIiImZmZmZmZd3d3ZmZmd3d3iIiImZmZiIiId3d3ZmZmVVVVZmZmZmZmZmZmiIiIiIiImZmZiIiIiIiId3d3d3d3d3d3d3d3ZmZmd3d3iIiIiIiIiIiIiIiIiIiId3d3VVVVZmZmZmZmZmZmVVVVZmZmiIiIqqqqu7u7u7u7u7u7u7u7zMzMu7u7qqqqiIiIZmZmd3d3iIiId3d3d3d3VVVVVVVVVVVVZmZmd3d3d3d3ZmZmZmZmVVVVd3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmVVVVd3d3d3d3mZmZmZmZmZmZiIiId3d3ZmZmiIiImZmZqqqqiIiIZmZmd3d3d3d3mZmZqqqqu7u7zMzMu7u7qqqqiIiId3d3d3d3d3d3d3d3ZmZmVVVVZmZmd3d3d3d3ZmZmZmZmZmZmiIiImZmZqqqqmZmZiIiId3d3ZmZmd3d3iIiIiIiImZmZiIiId3d3ZmZmiIiIiIiIiIiIZmZmVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmVVVVd3d3d3d3ZmZmVVVVREREVVVVVVVVVVVVZmZmiIiImZmZmZmZmZmZd3d3ZmZmiIiIu7u77u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////+7u7t3d3czMzMzMzLu7u8zMzN3d3e7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7u7u7u7u7t3d3czMzLu7u8zMzMzMzN3d3e7u7u7u7szMzLu7u8zMzN3d3d3d3czMzKqqqpmZmaqqqszMzN3d3d3d3d3d3czMzMzMzLu7u7u7u7u7u8zMzMzMzLu7u7u7u6qqqqqqqoiIiIiIiIiIiIiIiHd3d3d3d3d3d4iIiKqqqru7u8zMzN3d3e7u7t3d3d3d3czMzKqqqpmZmYiIiIiIiHd3d3d3d3d3d2ZmZnd3d3d3d4iIiHd3d3d3d3d3d3d3d2ZmZnd3d4iIiIiIiKqqqru7u7u7u8zMzN3d3czMzMzMzKqqqru7u6qqqqqqqpmZmYiIiIiIiHd3d3d3d3d3d3d3d2ZmZlVVVURERERERDMzM0RERERERFVVVVVVVVVVVWZmZmZmZmZmZlVVVWZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiHd3d4iIiJmZmZmZmbu7u8zMzMzMzN3d3czMzN3d3czMzLu7u7u7u7u7u8zMzN3d3bu7u7u7u8zMzLu7u5mZmXd3d2ZmZlVVVVVVVVVVVVVVVWZmZmZmZnd3d4iIiHd3d3d3d4iIiHd3d3d3d4iIiHd3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d2ZmZmZmZnd3d3d3d4iIiIiIiIiIiJmZmYiIiJmZmYiIiIiIiGZmZnd3d3d3d4iIiIiIiKqqqpmZmZmZmXd3d3d3d2ZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZlVVVWZmZnd3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d6qqqqqqqru7u6qqqqqqqpmZmZmZmZmZmaqqqru7u7u7u7u7u5mZmZmZmZmZmaqqqqqqqszMzMzMzLu7u7u7u7u7u5mZmZmZmYiIiIiIiIiIiIiIiHd3d3d3d2ZmZmZmZmZmZnd3d4iIiHd3d3d3d1VVVVVVVWZmZnd3d5mZmZmZmZmZmXd3d2ZmZnd3d5mZmaqqqru7u7u7u7u7u6qqqru7u6qqqqqqqqqqqqqqqqqqqqqqqru7u7u7u6qqqpmZmZmZmYiIiIiIiIiIiGZmZlVVVVVVVURERGZmZlVVVVVVVURERFVVVVVVVYiIiJmZmZmZmZmZmYiIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d4iIiIiIiGZmZmZmZnd3d4iIiIiIiIiIiGZmZmZmZmZmZlVVVVVVVWZmZnd3d3d3d4iIiIiIiHd3d3d3d3d3d3d3d3d3d2ZmZnd3d4iIiHd3d4iIiIiIiIiIiHd3d2ZmZlVVVWZmZnd3d2ZmZlVVVYiIiKqqqru7u7u7u7u7u7u7u7u7u7u7u6qqqpmZmYiIiHd3d3d3d3d3d2ZmZlVVVVVVVWZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZlVVVWZmZmZmZnd3d5mZmYiIiHd3d3d3d3d3d3d3d5mZmZmZmXd3d3d3d2ZmZnd3d5mZmZmZmaqqqru7u7u7u6qqqoiIiHd3d3d3d3d3d2ZmZmZmZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZnd3d6qqqqqqqpmZmYiIiHd3d2ZmZmZmZnd3d4iIiJmZmYiIiHd3d2ZmZnd3d4iIiIiIiGZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZoiIiHd3d3d3d2ZmZmZmZnd3d3d3d2ZmZlVVVURERERERERERGZmZnd3d4iIiJmZmYiIiHd3d2ZmZmZmZoiIiLu7u+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7d3d3d3d3d3d3MzMy7u7u7u7uZmZmIiIiIiIiZmZmqqqq7u7vMzMzd3d3d3d3u7u7u7u7u7u7u7u7u7u7d3d27u7uqqqqqqqq7u7u7u7vMzMzd3d2qqqqIiIiqqqqqqqqZmZmIiIhmZmZmZmaIiIi7u7vMzMzMzMzMzMzd3d3MzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3MzMy7u7uqqqqqqqqqqqqIiIiIiIhmZmZmZmZVVVVmZmZ3d3eZmZmZmZm7u7vMzMzd3d3d3d27u7u7u7uqqqqZmZmZmZmIiIiIiIh3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIh3d3d3d3dmZmZmZmZ3d3eIiIiIiIiqqqq7u7vMzMzMzMzMzMzMzMzMzMy7u7uZmZmZmZmIiIh3d3dmZmZVVVVmZmZVVVVVVVVVVVVVVVVEREREREQzMzMzMzNERERERERVVVVmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVmZmZ3d3dmZmZ3d3d3d3dmZmZ3d3d3d3d3d3eIiIiIiIiZmZm7u7u7u7vd3d3d3d3d3d3d3d27u7u7u7vMzMzd3d27u7uqqqqqqqrMzMy7u7uqqqqIiIh3d3d3d3dVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZ3d3d3d3d3d3eIiIh3d3dmZmZ3d3dmZmZ3d3d3d3eIiIiIiIiIiIiIiIh3d3d3d3eIiIh3d3eIiIiIiIiZmZmIiIiZmZmZmZmIiIh3d3d3d3d3d3eIiIiIiIiIiIiZmZmZmZmIiIhmZmZVVVVVVVVERERVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZ3d3d3d3eIiIiqqqqqqqqqqqqqqqqIiIiIiIiIiIiZmZm7u7u7u7u7u7uZmZmZmZmZmZmZmZmqqqqZmZmqqqqqqqqZmZmZmZmIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmaIiIh3d3d3d3dmZmZmZmZVVVVmZmZ3d3eIiIiIiIiIiIhmZmZmZmaIiIiZmZm7u7u7u7u7u7u7u7u7u7u7u7uqqqqqqqqqqqqqqqqqqqq7u7uqqqq7u7u7u7uZmZmIiIiIiIiIiIh3d3dmZmZmZmZVVVVVVVVVVVVmZmZVVVVERERVVVV3d3d3d3eIiIiIiIiZmZmqqqqqqqqqqqqZmZmZmZmZmZmZmZmIiIiIiIiIiIh3d3eIiIh3d3dmZmZmZmZmZmZ3d3d3d3eIiIhmZmZVVVVmZmZVVVVVVVVVVVV3d3eIiIiIiIiIiIh3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIiZmZmIiIh3d3dmZmZVVVVmZmZmZmZmZmZ3d3eZmZm7u7vMzMy7u7uqqqqZmZmqqqq7u7u7u7uZmZmIiIiIiIh3d3d3d3dmZmZVVVVVVVVmZmZmZmaIiIiIiIhmZmZVVVVmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZVVVV3d3eIiIiIiIiIiIiIiIh3d3d3d3eIiIiIiIh3d3dmZmZVVVVmZmaIiIiIiIiqqqqqqqq7u7uZmZmIiIh3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3eIiIhmZmZmZmZ3d3eZmZmqqqqqqqqIiIh3d3dVVVVVVVVmZmZ3d3eZmZmIiIhmZmZmZmZmZmaIiIiIiIhmZmZERERVVVVVVVVmZmZmZmZmZmZmZmZmZmaIiIh3d3d3d3dmZmZ3d3d3d3d3d3dmZmZVVVVERERERERERERVVVV3d3eIiIiIiIh3d3dmZmZVVVVmZmaIiIi7u7vd3d3///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////7u7u////////////////////7u7u////////////7u7u////////7u7u////////////////7u7u////////////////7u7u////////////7u7u////7u7u7u7u3d3d3d3dzMzMu7u7u7u7qqqqqqqqqqqqqqqqmZmZmZmZmZmZiIiImZmZqqqqzMzM3d3d3d3d7u7u7u7u7u7u3d3d3d3du7u7u7u7qqqqu7u7u7u7u7u7qqqqmZmZiIiIiIiId3d3d3d3ZmZmZmZmd3d3mZmZmZmZqqqqu7u7qqqqu7u7zMzMzMzM3d3d3d3d7u7u3d3d7u7u3d3d3d3d3d3dzMzMzMzMqqqqqqqqd3d3d3d3d3d3ZmZmZmZmd3d3d3d3d3d3iIiIiIiIqqqqqqqqu7u7zMzMu7u7u7u7qqqqqqqqmZmZiIiIiIiId3d3d3d3iIiIiIiIiIiIiIiIiIiId3d3d3d3VVVVVVVVZmZmZmZmiIiImZmZqqqqu7u7zMzMzMzMzMzMu7u7qqqqmZmZiIiIiIiIZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3iIiIiIiImZmZqqqqu7u7zMzMzMzMzMzMzMzM3d3d3d3dzMzMmZmZmZmZmZmZmZmZmZmZmZmZiIiImZmZiIiIZmZmVVVVVVVVREREREREREREVVVVZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiImZmZqqqqmZmZmZmZmZmZiIiId3d3iIiIiIiIiIiIiIiImZmZmZmZiIiIiIiIZmZmd3d3ZmZmd3d3iIiIiIiImZmZiIiId3d3d3d3VVVVVVVVVVVVVVVVZmZmZmZmd3d3ZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmZmZmZmZmd3d3d3d3iIiImZmZqqqqqqqqmZmZmZmZiIiIiIiId3d3iIiImZmZqqqqqqqqiIiIiIiId3d3d3d3d3d3d3d3iIiIiIiId3d3d3d3ZmZmd3d3d3d3ZmZmd3d3iIiId3d3ZmZmZmZmZmZmd3d3d3d3ZmZmd3d3d3d3ZmZmZmZmZmZmd3d3mZmZiIiId3d3d3d3d3d3mZmZu7u7u7u7zMzMu7u7u7u7qqqqmZmZqqqqqqqqqqqqqqqqqqqqu7u7u7u7u7u7mZmZiIiIiIiIiIiIiIiId3d3VVVVVVVVVVVVVVVVZmZmVVVVREREVVVVZmZmd3d3iIiImZmZqqqqqqqqu7u7u7u7u7u7u7u7qqqqmZmZmZmZiIiIiIiIiIiId3d3d3d3d3d3VVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmVVVVZmZmZmZmd3d3mZmZiIiIiIiId3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiId3d3ZmZmZmZmZmZmZmZmZmZmiIiImZmZu7u7u7u7u7u7qqqqmZmZqqqqu7u7u7u7qqqqmZmZd3d3d3d3d3d3d3d3VVVVVVVVZmZmd3d3d3d3d3d3ZmZmVVVVVVVVVVVVZmZmZmZmd3d3iIiId3d3iIiId3d3d3d3ZmZmZmZmZmZmZmZmd3d3iIiIiIiIiIiId3d3ZmZmd3d3iIiIiIiIZmZmZmZmVVVVZmZmd3d3iIiIiIiIqqqqmZmZmZmZd3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmd3d3d3d3ZmZmZmZmVVVVd3d3iIiImZmZiIiIiIiId3d3ZmZmREREZmZmd3d3iIiIiIiIZmZmVVVVZmZmiIiId3d3ZmZmVVVVREREVVVVZmZmZmZmZmZmZmZmd3d3iIiId3d3ZmZmZmZmZmZmd3d3ZmZmZmZmVVVVVVVVREREREREVVVVZmZmiIiImZmZiIiId3d3ZmZmd3d3d3d3mZmZ3d3d7u7u////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7t3d3d3d3czMzMzMzLu7u7u7u7u7u7u7u7u7u6qqqru7u6qqqqqqqpmZmZmZmaqqqqqqqru7u8zMzN3d3d3d3d3d3d3d3d3d3czMzLu7u8zMzLu7u7u7u7u7u6qqqpmZmZmZmZmZmZmZmZmZmYiIiIiIiHd3d4iIiJmZmaqqqpmZmaqqqqqqqru7u8zMzN3d3d3d3d3d3d3d3e7u7t3d3e7u7t3d3d3d3czMzMzMzLu7u5mZmYiIiHd3d3d3d4iIiHd3d3d3d4iIiHd3d3d3d3d3d3d3d5mZmZmZmbu7u7u7u8zMzLu7u7u7u6qqqpmZmYiIiIiIiJmZmYiIiIiIiIiIiIiIiHd3d4iIiGZmZmZmZlVVVVVVVVVVVWZmZnd3d5mZmZmZmaqqqru7u7u7u7u7u7u7u6qqqoiIiIiIiHd3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERDMzM0RERFVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZnd3d3d3d4iIiIiIiIiIiJmZmZmZmaqqqru7u8zMzMzMzMzMzMzMzMzMzLu7u7u7u5mZmYiIiHd3d3d3d4iIiJmZmaqqqpmZmYiIiGZmZlVVVURERERERERERFVVVURERFVVVVVVVWZmZmZmZnd3d3d3d4iIiJmZmZmZmaqqqru7u7u7u6qqqru7u6qqqqqqqpmZmZmZmYiIiIiIiIiIiIiIiIiIiJmZmYiIiIiIiGZmZnd3d2ZmZnd3d4iIiIiIiIiIiIiIiIiIiHd3d2ZmZlVVVVVVVURERGZmZmZmZmZmZnd3d2ZmZnd3d2ZmZmZmZlVVVWZmZnd3d2ZmZlVVVWZmZmZmZmZmZnd3d3d3d4iIiIiIiIiIiIiIiJmZmaqqqqqqqpmZmYiIiIiIiIiIiHd3d4iIiJmZmZmZmYiIiGZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d2ZmZlVVVWZmZnd3d5mZmYiIiHd3d2ZmZnd3d5mZmbu7u7u7u7u7u6qqqqqqqpmZmZmZmaqqqqqqqqqqqqqqqqqqqru7u6qqqpmZmYiIiIiIiIiIiIiIiIiIiGZmZlVVVURERERERFVVVVVVVURERERERFVVVXd3d3d3d5mZmaqqqqqqqru7u7u7u8zMzMzMzLu7u5mZmZmZmZmZmYiIiIiIiHd3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZlVVVWZmZmZmZlVVVVVVVWZmZmZmZoiIiJmZmYiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d4iIiJmZmYiIiHd3d2ZmZmZmZmZmZmZmZnd3d2ZmZoiIiKqqqru7u7u7u6qqqpmZmZmZmZmZmbu7u6qqqpmZmYiIiIiIiHd3d3d3d2ZmZmZmZlVVVWZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZnd3d4iIiIiIiIiIiHd3d2ZmZmZmZmZmZmZmZnd3d3d3d4iIiIiIiHd3d2ZmZmZmZmZmZnd3d3d3d2ZmZlVVVVVVVWZmZnd3d4iIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d4iIiHd3d2ZmZmZmZmZmZnd3d2ZmZmZmZlVVVWZmZmZmZmZmZoiIiIiIiHd3d3d3d2ZmZlVVVVVVVXd3d5mZmYiIiGZmZmZmZmZmZoiIiHd3d2ZmZkRERFVVVVVVVWZmZnd3d2ZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZmZmZnd3d2ZmZlVVVURERFVVVURERFVVVWZmZnd3d5mZmYiIiHd3d2ZmZmZmZnd3d4iIiN3d3f///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP//AAD//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7u7u7t3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u7u7u6qqqru7u6qqqru7u7u7u7u7u7u7u7u7u7u7u7u7u8zMzLu7u8zMzMzMzLu7u7u7u7u7u6qqqqqqqqqqqqqqqru7u7u7u6qqqqqqqqqqqqqqqpmZmaqqqqqqqru7u7u7u8zMzMzMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzLu7u7u7u6qqqqqqqqqqqpmZmZmZmZmZmYiIiIiIiHd3d4iIiHd3d3d3d3d3d4iIiJmZmZmZmbu7u7u7u7u7u7u7u6qqqqqqqpmZmZmZmYiIiIiIiIiIiHd3d2ZmZnd3d3d3d3d3d2ZmZmZmZlVVVVVVVVVVVWZmZnd3d3d3d4iIiJmZmZmZmaqqqru7u7u7u6qqqoiIiIiIiHd3d3d3d2ZmZmZmZlVVVVVVVWZmZlVVVWZmZlVVVVVVVVVVVURERERERERERERERFVVVVVVVWZmZnd3d2ZmZnd3d2ZmZmZmZmZmZnd3d3d3d3d3d4iIiIiIiIiIiJmZmZmZmZmZmZmZmaqqqqqqqru7u8zMzN3d3czMzMzMzLu7u7u7u5mZmYiIiHd3d3d3d3d3d3d3d5mZmZmZmZmZmYiIiGZmZlVVVURERERERFVVVVVVVXd3d2ZmZnd3d4iIiIiIiJmZmbu7u8zMzLu7u8zMzMzMzMzMzMzMzMzMzLu7u7u7u6qqqpmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d2ZmZnd3d3d3d4iIiIiIiIiIiIiIiIiIiHd3d2ZmZlVVVURERFVVVVVVVWZmZmZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZoiIiIiIiIiIiIiIiIiIiJmZmZmZmaqqqqqqqpmZmZmZmZmZmXd3d4iIiIiIiIiIiIiIiGZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d3d3d3d3d2ZmZnd3d2ZmZmZmZmZmZlVVVWZmZnd3d3d3d3d3d3d3d1VVVVVVVWZmZnd3d4iIiIiIiHd3d2ZmZnd3d3d3d5mZmaqqqru7u6qqqqqqqqqqqqqqqqqqqpmZmZmZmbu7u6qqqpmZmZmZmYiIiHd3d3d3d3d3d5mZmaqqqoiIiGZmZkRERERERERERERERERERFVVVVVVVWZmZoiIiJmZmaqqqszMzMzMzMzMzMzMzMzMzMzMzKqqqqqqqpmZmZmZmXd3d3d3d3d3d3d3d1VVVWZmZmZmZmZmZnd3d2ZmZlVVVVVVVVVVVVVVVXd3d2ZmZlVVVVVVVXd3d4iIiHd3d3d3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d4iIiJmZmXd3d2ZmZmZmZmZmZnd3d3d3d2ZmZoiIiJmZmaqqqru7u6qqqqqqqpmZmZmZmaqqqqqqqqqqqoiIiIiIiIiIiHd3d3d3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVXd3d4iIiIiIiIiIiHd3d3d3d2ZmZnd3d2ZmZnd3d3d3d4iIiJmZmZmZmXd3d2ZmZlVVVWZmZmZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZoiIiHd3d3d3d3d3d3d3d3d3d4iIiHd3d2ZmZmZmZlVVVWZmZmZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZnd3d3d3d3d3d2ZmZlVVVVVVVXd3d4iIiIiIiHd3d1VVVWZmZoiIiHd3d2ZmZlVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d4iIiHd3d3d3d3d3d3d3d2ZmZmZmZlVVVURERFVVVURERFVVVVVVVXd3d4iIiKqqqoiIiFVVVVVVVWZmZoiIiMzMzP///////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7d3d3d3d3MzMzMzMzd3d3d3d3d3d3d3d3MzMzMzMzMzMy7u7u7u7u7u7uqqqqqqqq7u7uqqqqqqqq7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7vMzMy7u7u7u7vMzMy7u7u7u7u7u7u7u7uqqqq7u7u7u7u7u7u7u7vMzMzMzMzMzMzMzMzMzMzMzMzMzMy7u7u7u7uqqqq7u7u7u7u7u7u7u7u7u7uqqqqqqqqqqqqZmZmZmZmZmZmIiIiIiIh3d3d3d3d3d3d3d3eIiIiIiIiZmZmZmZm7u7u7u7uqqqqZmZmZmZmIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZ3d3eIiIiqqqqqqqqqqqqqqqqZmZmIiIh3d3dmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVERERERERERERERERVVVVVVVVmZmZ3d3d3d3d3d3eIiIiZmZmZmZmZmZmZmZmZmZmZmZmqqqqqqqqZmZmqqqqqqqqqqqqqqqq7u7u7u7vMzMzMzMzMzMzMzMyqqqqZmZmIiIh3d3dmZmZ3d3d3d3eZmZmZmZmZmZmIiIh3d3dVVVVmZmZmZmZmZmZ3d3d3d3eIiIiZmZmqqqq7u7vMzMzMzMzMzMzd3d3MzMzMzMzMzMzMzMy7u7vMzMyqqqqZmZmZmZl3d3d3d3d3d3eIiIiIiIiIiIiZmZl3d3dmZmZmZmZmZmZ3d3d3d3eIiIiIiIiIiIh3d3d3d3dVVVVVVVVVVVVVVVVVVVVERERVVVVmZmZVVVVVVVVmZmZmZmZVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3eIiIiZmZmZmZmZmZmZmZmZmZmqqqq7u7uqqqqZmZmIiIh3d3d3d3d3d3eIiIh3d3dmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3dmZmZVVVVVVVV3d3d3d3d3d3d3d3dmZmZmZmZ3d3eIiIiqqqq7u7uqqqq7u7uqqqqZmZmZmZmqqqqqqqqZmZmZmZmIiIiIiIiIiIh3d3d3d3eIiIiqqqqZmZmIiIhmZmZERERERERERERVVVVERERVVVVVVVV3d3eZmZmqqqq7u7vMzMzMzMzd3d3MzMzMzMzMzMy7u7u7u7uqqqqZmZmIiIh3d3d3d3d3d3dmZmZmZmZVVVVmZmZmZmZVVVVERERVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3eIiIiqqqqIiIhmZmaIiIiZmZmqqqp3d3dmZmZmZmZmZmZmZmZ3d3dmZmZ3d3eIiIiqqqrMzMy7u7vMzMyZmZmZmZmZmZm7u7uqqqqIiIh3d3d3d3d3d3dmZmZmZmZmZmZVVVVVVVVERERERERVVVVERERVVVVVVVVmZmZ3d3d3d3eIiIh3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3eZmZmqqqqIiIhmZmZmZmZVVVVVVVVVVVVVVVVERERERERVVVVVVVV3d3eIiIiIiIh3d3dmZmZmZmZmZmZ3d3eIiIh3d3d3d3dmZmZmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmaIiIiIiIh3d3dmZmZERERVVVWZmZmqqqqIiIh3d3dVVVVmZmaIiIh3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZ3d3d3d3eIiIiIiIiIiIiIiIh3d3dmZmZmZmZVVVVERERERERERERVVVVVVVVmZmaZmZmZmZl3d3dVVVVVVVVmZmaZmZnd3d3////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////7u7u7u7u7u7u3d3d3d3d3d3d7u7u7u7u7u7u7u7u3d3d3d3dzMzMzMzMu7u7u7u7qqqqmZmZmZmZiIiImZmZmZmZqqqqqqqqqqqqu7u7u7u7u7u7zMzMzMzMzMzMzMzM3d3dzMzMzMzMzMzMu7u7qqqqmZmZmZmZmZmZmZmZmZmZmZmZqqqqmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZqqqqqqqqqqqqqqqqu7u7u7u7u7u7qqqqqqqqmZmZmZmZiIiIiIiId3d3d3d3d3d3ZmZmZmZmd3d3d3d3mZmZmZmZqqqqqqqqmZmZmZmZmZmZiIiIiIiId3d3iIiIiIiId3d3d3d3ZmZmVVVVZmZmVVVVVVVVREREVVVVREREREREVVVVZmZmd3d3iIiImZmZmZmZmZmZmZmZiIiId3d3ZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmd3d3d3d3iIiIqqqqqqqqqqqqqqqqqqqqmZmZmZmZqqqqqqqqmZmZqqqqqqqqqqqqqqqqqqqqqqqqu7u7zMzMzMzMzMzMu7u7u7u7qqqqiIiId3d3ZmZmVVVVd3d3d3d3mZmZiIiIiIiIiIiIZmZmZmZmZmZmd3d3iIiIqqqqu7u7u7u7u7u7zMzMzMzM3d3dzMzMzMzMzMzMzMzMu7u7u7u7zMzMu7u7qqqqmZmZiIiIiIiId3d3d3d3d3d3mZmZiIiIiIiIZmZmZmZmZmZmd3d3iIiId3d3iIiIiIiIiIiIiIiId3d3ZmZmVVVVVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmd3d3d3d3iIiIiIiImZmZmZmZmZmZmZmZqqqqqqqqu7u7u7u7mZmZmZmZiIiId3d3ZmZmZmZmd3d3ZmZmZmZmVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmZmZmd3d3iIiImZmZmZmZiIiIZmZmVVVVd3d3d3d3d3d3d3d3ZmZmVVVVZmZmd3d3mZmZqqqqqqqqqqqqmZmZmZmZmZmZmZmZmZmZiIiImZmZd3d3d3d3d3d3d3d3d3d3d3d3mZmZmZmZd3d3VVVVREREREREREREREREVVVVZmZmZmZmiIiIqqqqu7u7u7u7u7u7u7u7zMzMzMzM3d3dzMzMu7u7u7u7u7u7mZmZiIiId3d3d3d3d3d3ZmZmVVVVVVVVVVVVVVVVVVVVREREREREVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVd3d3iIiIiIiIiIiId3d3d3d3iIiIu7u7qqqqd3d3VVVVVVVVZmZmd3d3ZmZmVVVVd3d3mZmZqqqqu7u7zMzMu7u7qqqqmZmZmZmZqqqqu7u7mZmZd3d3d3d3d3d3iIiId3d3ZmZmVVVVVVVVREREREREREREVVVVVVVVVVVVd3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3iIiIqqqqmZmZmZmZiIiIZmZmREREREREVVVVREREREREREREVVVVZmZmiIiId3d3d3d3d3d3ZmZmVVVVZmZmd3d3d3d3d3d3ZmZmZmZmVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmd3d3iIiId3d3ZmZmVVVVZmZmiIiIqqqqmZmZiIiIZmZmVVVVZmZmiIiIZmZmREREREREREREZmZmZmZmVVVVVVVVd3d3iIiImZmZiIiIiIiIiIiId3d3VVVVZmZmVVVVREREREREREREREREVVVVVVVVZmZmiIiIiIiIZmZmVVVVVVVVVVVVmZmZ3d3d////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7v///+7u7v///////////////////////////////////////+7u7v///////////////////+7u7v///////////+7u7v///////////////////////////////////////////////////////////////////+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3czMzMzMzKqqqpmZmYiIiHd3d3d3d3d3d4iIiKqqqqqqqru7u8zMzMzMzLu7u8zMzMzMzMzMzMzMzMzMzLu7u7u7u6qqqpmZmYiIiIiIiHd3d3d3d3d3d3d3d3d3d2ZmZmZmZnd3d3d3d3d3d4iIiIiIiIiIiIiIiJmZmYiIiJmZmZmZmaqqqqqqqpmZmZmZmYiIiIiIiIiIiHd3d3d3d3d3d2ZmZmZmZlVVVVVVVWZmZmZmZnd3d4iIiJmZmZmZmZmZmZmZmYiIiJmZmYiIiIiIiIiIiHd3d2ZmZmZmZlVVVWZmZlVVVVVVVVVVVVVVVURERFVVVURERFVVVVVVVXd3d3d3d4iIiJmZmaqqqoiIiHd3d3d3d3d3d2ZmZmZmZnd3d2ZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d2ZmZoiIiJmZmZmZmZmZmaqqqqqqqqqqqqqqqqqqqpmZmaqqqqqqqqqqqpmZmZmZmaqqqpmZmaqqqqqqqqqqqqqqqru7u8zMzMzMzMzMzKqqqpmZmZmZmYiIiFVVVVVVVWZmZnd3d4iIiJmZmZmZmYiIiIiIiHd3d4iIiJmZmZmZmaqqqru7u7u7u7u7u7u7u8zMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u7u7u6qqqqqqqpmZmYiIiHd3d2ZmZnd3d4iIiIiIiIiIiHd3d2ZmZmZmZlVVVWZmZnd3d3d3d4iIiIiIiIiIiIiIiGZmZmZmZlVVVURERERERFVVVURERFVVVVVVVWZmZmZmZmZmZmZmZnd3d3d3d4iIiIiIiJmZmZmZmZmZmZmZmbu7u6qqqqqqqqqqqru7u7u7u6qqqpmZmZmZmYiIiHd3d2ZmZmZmZmZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVWZmZlVVVWZmZmZmZlVVVWZmZmZmZmZmZmZmZnd3d4iIiHd3d3d3d3d3d1VVVVVVVWZmZnd3d3d3d2ZmZmZmZlVVVWZmZmZmZoiIiIiIiJmZmZmZmYiIiIiIiJmZmYiIiIiIiIiIiHd3d2ZmZmZmZmZmZnd3d3d3d3d3d4iIiIiIiGZmZlVVVURERERERERERFVVVVVVVXd3d3d3d5mZmaqqqru7u8zMzLu7u8zMzMzMzMzMzMzMzMzMzMzMzMzMzKqqqpmZmYiIiGZmZmZmZnd3d2ZmZmZmZlVVVVVVVURERERERERERERERFVVVWZmZmZmZnd3d2ZmZlVVVVVVVVVVVVVVVWZmZnd3d4iIiHd3d3d3d3d3d3d3d5mZmbu7u3d3d2ZmZlVVVVVVVWZmZlVVVVVVVVVVVWZmZoiIiKqqqru7u6qqqqqqqpmZmZmZmaqqqru7u5mZmYiIiGZmZnd3d4iIiHd3d2ZmZmZmZlVVVVVVVURERERERERERERERFVVVWZmZlVVVVVVVWZmZmZmZmZmZnd3d3d3d4iIiHd3d3d3d4iIiJmZmZmZmaqqqoiIiHd3d1VVVURERDMzM0RERERERERERFVVVWZmZnd3d3d3d2ZmZmZmZnd3d3d3d2ZmZmZmZmZmZnd3d3d3d2ZmZmZmZlVVVWZmZmZmZmZmZkRERERERFVVVVVVVWZmZnd3d3d3d2ZmZlVVVXd3d5mZmZmZmYiIiJmZmZmZmWZmZkRERFVVVVVVVURERDMzMzMzM1VVVXd3d2ZmZmZmZmZmZnd3d3d3d4iIiIiIiIiIiHd3d3d3d3d3d2ZmZlVVVVVVVVVVVURERFVVVVVVVWZmZnd3d4iIiIiIiHd3d2ZmZmZmZmZmZqqqqu7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3d3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7////u7u7u7u7u7u7u7u7d3d3d3d3d3d3u7u7u7u7////////u7u7////////////u7u7////////d3d3MzMzu7u7////////////////////////////////////////////////////////////u7u7////u7u7////u7u7////u7u7u7u7u7u7d3d3MzMy7u7uqqqqIiIhmZmZmZmZ3d3d3d3eIiIiqqqq7u7u7u7vMzMzMzMzMzMzMzMzMzMy7u7uqqqqZmZmIiIiZmZl3d3eIiIh3d3eIiIiIiIh3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIh3d3d3d3dmZmZmZmZmZmZVVVVmZmZmZmZVVVVVVVVVVVVERERERERVVVVmZmZmZmZ3d3eIiIiIiIiZmZmZmZmZmZmIiIiIiIiIiIh3d3dmZmZmZmZmZmZVVVVVVVVmZmZVVVVVVVVERERVVVVVVVVERERVVVVVVVVmZmZ3d3eIiIiZmZmZmZmIiIiIiIh3d3d3d3eIiIh3d3dmZmZmZmZmZmZmZmZmZmZ3d3d3d3eIiIiIiIiIiIiIiIiIiIiZmZmIiIiZmZmIiIiZmZmqqqqqqqqqqqq7u7uqqqq7u7u7u7uqqqqqqqqqqqqZmZmZmZmZmZmIiIiZmZmZmZmqqqqZmZmqqqqqqqq7u7u7u7uqqqqZmZl3d3dmZmZVVVVmZmZmZmaIiIiZmZmZmZmqqqqZmZmZmZmZmZmZmZmIiIiZmZmqqqq7u7u7u7u7u7vMzMzMzMzMzMzMzMy7u7u7u7u7u7uqqqq7u7uqqqqqqqqIiIh3d3dmZmZmZmZ3d3d3d3eIiIiIiIh3d3dmZmZVVVVmZmZmZmZ3d3d3d3eIiIiZmZmIiIiIiIh3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3eZmZmIiIiZmZmqqqqZmZmqqqqqqqqqqqqqqqqqqqqqqqqqqqq7u7u7u7u7u7uqqqqZmZmZmZmIiIh3d3dVVVVmZmZVVVVVVVVVVVVERERERERVVVVmZmZ3d3dmZmZVVVVERERVVVVERERVVVVVVVVVVVVmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZERERVVVVVVVVmZmZ3d3d3d3dVVVVVVVVERERVVVVVVVV3d3d3d3eIiIiIiIh3d3d3d3d3d3d3d3dmZmZ3d3dmZmZmZmZmZmZ3d3d3d3d3d3eIiIiIiIh3d3dmZmZVVVVVVVVERERERERVVVVmZmZ3d3d3d3eIiIiZmZmqqqrMzMy7u7u7u7u7u7u7u7vMzMzd3d3d3d3d3d27u7uZmZl3d3dmZmZ3d3d3d3d3d3dVVVVVVVVVVVVEREQzMzMzMzNERERERERVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3dmZmZ3d3d3d3eIiIiIiIhVVVVERERVVVVVVVVVVVVVVVVVVVVVVVV3d3eZmZmZmZmZmZmqqqqqqqqZmZmZmZmqqqqZmZmIiIh3d3dVVVVVVVVmZmZ3d3dmZmZmZmZEREQzMzMzMzMzMzNERERERERERERERERVVVVERERVVVVmZmZmZmZ3d3d3d3d3d3eZmZmZmZmIiIiIiIh3d3dmZmZVVVVEREREREQzMzNEREQzMzNERERVVVVVVVVVVVVVVVVERERmZmaIiIiIiIhmZmZmZmZmZmZmZmaIiIiIiIhmZmZVVVVmZmZmZmZVVVVERERERERVVVVmZmZmZmZVVVVVVVVERERVVVV3d3d3d3d3d3eZmZmqqqqZmZlmZmZEREREREREREQzMzMiIiIzMzNERERmZmZ3d3dmZmZmZmZmZmZ3d3d3d3eIiIiIiIiZmZmIiIh3d3dVVVVVVVVVVVVERERVVVVERERVVVV3d3d3d3eZmZmqqqp3d3dmZmZVVVVmZmaqqqru7u7////u7u7////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u////7u7u7u7u3d3d3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzMzMzMzMzMu7u7qqqqzMzM3d3d3d3d7u7u7u7u7u7u7u7u////7u7u////////////////////////////////////7u7u////////7u7u7u7u7u7u3d3d3d3dzMzMzMzMu7u7mZmZiIiIZmZmZmZmZmZmVVVVZmZmiIiIiIiIqqqqu7u7u7u7zMzMzMzMu7u7u7u7qqqqmZmZiIiIiIiIiIiIiIiImZmZmZmZmZmZmZmZiIiId3d3d3d3d3d3ZmZmVVVVVVVVVVVVZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVZmZmVVVVVVVVVVVVREREREREVVVVREREVVVVZmZmiIiIiIiIiIiImZmZiIiIqqqqmZmZd3d3iIiIZmZmZmZmZmZmVVVVZmZmVVVVREREVVVVREREVVVVREREREREVVVVREREVVVVZmZmd3d3iIiImZmZmZmZiIiIiIiIiIiId3d3d3d3ZmZmZmZmZmZmZmZmd3d3iIiIiIiImZmZiIiImZmZiIiIiIiIiIiIiIiImZmZmZmZqqqqqqqqqqqqzMzMu7u7u7u7u7u7qqqqqqqqqqqqmZmZmZmZmZmZiIiImZmZiIiIiIiIiIiId3d3mZmZqqqqqqqqqqqqqqqqmZmZd3d3d3d3ZmZmZmZmd3d3d3d3iIiIqqqqu7u7u7u7mZmZmZmZmZmZmZmZmZmZqqqqqqqqu7u7u7u7u7u7zMzMzMzMu7u7u7u7u7u7qqqqqqqqqqqqmZmZiIiId3d3VVVVVVVVZmZmZmZmd3d3iIiId3d3ZmZmVVVVVVVVZmZmZmZmd3d3d3d3iIiIiIiImZmZiIiId3d3VVVVVVVVVVVVVVVVZmZmd3d3ZmZmd3d3iIiImZmZqqqqqqqqmZmZqqqqqqqqqqqqmZmZqqqqmZmZqqqqqqqqmZmZqqqqu7u7u7u7qqqqqqqqmZmZmZmZiIiId3d3VVVVVVVVREREREREVVVVREREREREVVVVVVVVVVVVVVVVREREREREVVVVVVVVVVVVVVVVZmZmd3d3ZmZmZmZmZmZmd3d3ZmZmZmZmVVVVVVVVVVVVd3d3ZmZmZmZmVVVVREREREREREREVVVVZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmd3d3d3d3d3d3d3d3iIiImZmZd3d3VVVVREREREREREREVVVVVVVVVVVVZmZmd3d3mZmZqqqqqqqqqqqqqqqqu7u7qqqqu7u7zMzM3d3d3d3du7u7iIiIZmZmd3d3mZmZiIiIVVVVVVVVVVVVREREMzMzMzMzMzMzREREREREREREREREVVVVVVVVVVVVZmZmVVVVVVVVVVVVZmZmZmZmd3d3iIiIZmZmZmZmiIiIiIiIVVVVVVVVREREREREREREREREREREREREREREVVVVZmZmd3d3iIiIiIiImZmZiIiIiIiIiIiImZmZmZmZZmZmREREVVVVZmZmVVVVREREREREMzMzREREMzMzMzMzREREREREREREREREREREREREVVVVVVVVVVVVZmZmZmZmiIiIiIiIZmZmVVVVVVVVZmZmVVVVVVVVVVVVREREREREREREMzMzMzMzREREREREREREMzMzVVVVZmZmd3d3ZmZmVVVVZmZmVVVVd3d3iIiIZmZmREREREREVVVVREREREREREREVVVVZmZmZmZmVVVVREREMzMzREREREREd3d3d3d3ZmZmiIiImZmZd3d3REREREREMzMzMzMzIiIiIiIiIiIiVVVVZmZmZmZmVVVVVVVVd3d3d3d3d3d3d3d3iIiImZmZiIiIZmZmVVVVVVVVVVVVREREVVVVZmZmVVVVd3d3iIiImZmZmZmZiIiIZmZmVVVVd3d3u7u77u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////+7u7v///////////////+7u7v///////////////////////////////////////////////////////+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7t3d3e7u7t3d3czMzMzMzMzMzLu7u7u7u7u7u7u7u6qqqqqqqpmZmaqqqszMzMzMzMzMzMzMzN3d3d3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7v///+7u7v///////////+7u7u7u7t3d3d3d3czMzMzMzLu7u6qqqpmZmZmZmYiIiHd3d2ZmZmZmZlVVVVVVVVVVVWZmZmZmZnd3d5mZmZmZmbu7u8zMzLu7u7u7u6qqqpmZmZmZmYiIiJmZmZmZmaqqqpmZmZmZmZmZmZmZmZmZmYiIiIiIiGZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVWZmZnd3d4iIiJmZmaqqqpmZmZmZmYiIiIiIiGZmZmZmZnd3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERFVVVVVVVWZmZoiIiIiIiJmZmZmZmYiIiHd3d3d3d2ZmZnd3d3d3d3d3d3d3d4iIiHd3d5mZmYiIiIiIiJmZmZmZmZmZmZmZmZmZmZmZmZmZmaqqqqqqqru7u6qqqru7u7u7u7u7u6qqqqqqqqqqqpmZmYiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d4iIiJmZmaqqqqqqqpmZmYiIiJmZmYiIiGZmZmZmZnd3d4iIiJmZmaqqqru7u7u7u6qqqpmZmZmZmZmZmZmZmZmZmbu7u6qqqru7u7u7u7u7u7u7u6qqqqqqqqqqqpmZmZmZmYiIiHd3d3d3d2ZmZlVVVVVVVWZmZnd3d3d3d3d3d2ZmZmZmZlVVVVVVVVVVVWZmZnd3d3d3d4iIiIiIiIiIiHd3d2ZmZlVVVWZmZmZmZnd3d3d3d4iIiJmZmaqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqpmZmaqqqqqqqpmZmaqqqqqqqqqqqqqqqqqqqpmZmYiIiHd3d1VVVURERFVVVURERERERERERFVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d2ZmZlVVVVVVVVVVVVVVVWZmZlVVVURERERERDMzM0RERERERFVVVWZmZmZmZmZmZnd3d3d3d2ZmZnd3d2ZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZnd3d6qqqqqqqmZmZkRERERERERERFVVVVVVVVVVVVVVVVVVVWZmZnd3d5mZmZmZmZmZmZmZmZmZmZmZmaqqqszMzN3d3bu7u4iIiHd3d2ZmZnd3d3d3d2ZmZlVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERFVVVWZmZlVVVURERFVVVWZmZnd3d1VVVVVVVWZmZmZmZkRERERERERERERERERERDMzM0RERERERERERDMzM0RERFVVVVVVVWZmZmZmZmZmZnd3d3d3d4iIiJmZmXd3d1VVVURERFVVVVVVVURERERERDMzM0RERDMzMzMzMzMzM0RERERERERERERERERERDMzM0RERERERERERERERFVVVVVVVURERFVVVURERFVVVVVVVVVVVVVVVURERERERDMzM0RERDMzMzMzMyIiIjMzMzMzMzMzM0RERGZmZlVVVURERERERFVVVVVVVWZmZlVVVVVVVVVVVURERERERDMzM0RERERERERERERERERERERERERERERERERERGZmZnd3d2ZmZmZmZnd3d4iIiHd3d1VVVURERDMzMyIiIiIiIiIiIjMzMzMzM0RERFVVVVVVVVVVVXd3d4iIiHd3d3d3d3d3d4iIiHd3d1VVVVVVVURERFVVVVVVVWZmZmZmZlVVVXd3d5mZmZmZmZmZmXd3d2ZmZlVVVXd3d8zMzO7u7u7u7v///////////+7u7v///////////+7u7v///////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////+7u7v///////////////////////////////////////////////////////////////////////////////+7u7v///////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////u7u7u7u7u7u7////u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3MzMzMzMzMzMy7u7u7u7u7u7vMzMzMzMzMzMzMzMzd3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7////u7u7////u7u7d3d3d3d27u7u7u7u7u7uqqqqqqqqZmZmZmZmIiIiIiIh3d3eIiIh3d3d3d3dmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZ3d3eIiIiqqqqZmZmqqqqqqqqqqqqZmZmIiIiqqqqZmZmZmZmZmZmqqqqqqqqZmZmZmZmIiIiIiIiIiIh3d3dmZmZmZmZVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERVVVVmZmZmZmaIiIiZmZmZmZmZmZmZmZmIiIiIiIiIiIh3d3d3d3dmZmZVVVVVVVVVVVVVVVVERERERERERERERERERERERERVVVVVVVVmZmZ3d3eIiIiqqqqqqqqZmZmZmZmIiIiIiIiIiIiZmZmZmZmIiIiIiIh3d3eIiIiIiIiZmZmZmZmZmZmqqqqZmZmZmZmZmZmZmZmZmZmZmZmqqqqqqqq7u7u7u7uqqqqqqqqZmZmIiIiIiIh3d3dmZmZmZmZVVVVVVVVVVVVVVVVmZmZ3d3eIiIiIiIiZmZmqqqqZmZmZmZmIiIiIiIiZmZmIiIiIiIiqqqq7u7u7u7u7u7u7u7uqqqqZmZmZmZmIiIiZmZmZmZmZmZmqqqqZmZmZmZmqqqqqqqqZmZmIiIh3d3d3d3dmZmZ3d3dmZmZVVVVVVVVERERVVVVmZmZ3d3d3d3dmZmZVVVVVVVVVVVVVVVVmZmZmZmZ3d3eIiIiZmZmIiIh3d3dmZmZmZmZmZmZ3d3d3d3eZmZmqqqqqqqqqqqqqqqqqqqqqqqq7u7u7u7uqqqq7u7u7u7uqqqqqqqqZmZmZmZmZmZmZmZmZmZmqqqqZmZmZmZmIiIiIiIhmZmZVVVVERERERERERERERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3dmZmZVVVVERERVVVVERERmZmZVVVVERERERERERERERERERERERERVVVVmZmZmZmZ3d3dmZmZmZmZmZmZVVVVmZmZVVVVmZmZmZmZmZmZ3d3d3d3eZmZmqqqp3d3dVVVUzMzNERERERERERERERERERERVVVVERERERERmZmZmZmZmZmaIiIiIiIh3d3eIiIiIiIiZmZm7u7uqqqp3d3dmZmZVVVVmZmZmZmZVVVVEREQzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERERERERERERERVVVVVVVVEREREREREREQzMzNEREQzMzMzMzMzMzMzMzNEREQzMzNEREREREQzMzMzMzMzMzNERERERERERERVVVVmZmZmZmZVVVVVVVVEREREREREREREREQzMzNEREREREREREREREQzMzMzMzNEREQzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNERERERERVVVVVVVVEREREREREREREREQzMzMzMzNEREQzMzMzMzNEREREREQzMzMzMzMzMzNERERVVVUzMzNVVVV3d3eIiIiIiIhEREQzMzNEREQiIiIiIiIiIiIiIiIiIiIzMzNERERERERmZmZ3d3eIiIiIiIhmZmZmZmaIiIhmZmZVVVVERERERERVVVVmZmZmZmZVVVVmZmZ3d3eIiIiZmZmZmZlmZmZVVVVVVVWIiIjd3d3////////////////////////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////7u7u////////////7u7u////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u3d3d7u7u7u7u3d3dzMzM3d3d3d3dzMzMzMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u3d3dzMzMu7u7mZmZmZmZmZmZiIiImZmZiIiIiIiIiIiId3d3d3d3d3d3d3d3ZmZmd3d3d3d3ZmZmd3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3mZmZmZmZmZmZqqqqqqqqmZmZmZmZmZmZmZmZqqqqmZmZmZmZmZmZmZmZmZmZd3d3d3d3d3d3ZmZmZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREVVVVREREVVVVZmZmZmZmVVVVREREVVVVVVVVREREVVVVREREREREVVVVVVVVZmZmd3d3iIiImZmZqqqqmZmZmZmZiIiIiIiId3d3ZmZmZmZmVVVVVVVVVVVVREREREREREREREREREREREREREREREREVVVVVVVVd3d3iIiImZmZqqqqmZmZmZmZqqqqu7u7u7u7qqqqmZmZmZmZiIiIiIiIiIiImZmZmZmZqqqqmZmZmZmZiIiIiIiIiIiIiIiIiIiIiIiImZmZmZmZmZmZiIiIiIiId3d3ZmZmZmZmVVVVREREVVVVREREREREVVVVREREVVVVVVVVZmZmd3d3iIiIiIiIqqqqqqqqmZmZqqqqmZmZiIiIiIiIiIiImZmZqqqqqqqqu7u7u7u7qqqqmZmZiIiIiIiIiIiId3d3iIiIiIiIiIiImZmZiIiIiIiId3d3d3d3d3d3d3d3d3d3ZmZmZmZmVVVVVVVVVVVVZmZmd3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVd3d3d3d3iIiImZmZiIiIiIiId3d3ZmZmZmZmZmZmiIiImZmZmZmZmZmZu7u7qqqqu7u7u7u7u7u7u7u7u7u7u7u7qqqqqqqqqqqqmZmZqqqqmZmZmZmZqqqqqqqqqqqqmZmZmZmZiIiId3d3VVVVREREREREREREMzMzMzMzMzMzMzMzREREVVVVREREVVVVZmZmVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmd3d3d3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmiIiIiIiIZmZmZmZmd3d3ZmZmREREMzMzMzMzREREREREREREREREREREMzMzMzMzMzMzREREREREVVVVVVVVZmZmVVVVZmZmiIiImZmZd3d3ZmZmVVVVVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzREREMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzREREMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiERERIiIiIiIiMzMzMzMzMzMzMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzREREVVVVZmZmVVVVREREREREMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzVVVVZmZmd3d3iIiId3d3ZmZmZmZmVVVVREREREREREREREREVVVVVVVVZmZmVVVVZmZmiIiImZmZqqqqd3d3VVVVVVVVVVVViIiIzMzM////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7v///+7u7u7u7u7u7u7u7u7u7v///////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7u7u7v///+7u7u7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3czMzMzMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3czMzLu7u5mZmYiIiHd3d4iIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZnd3d2ZmZnd3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d5mZmZmZmaqqqpmZmYiIiJmZmZmZmaqqqqqqqqqqqqqqqpmZmZmZmZmZmYiIiIiIiHd3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVURERERERDMzM0RERERERERERFVVVVVVVVVVVURERFVVVVVVVVVVVURERFVVVVVVVURERFVVVVVVVWZmZnd3d4iIiIiIiIiIiKqqqqqqqpmZmYiIiIiIiHd3d2ZmZmZmZlVVVVVVVURERERERERERERERERERFVVVURERFVVVVVVVVVVVWZmZoiIiIiIiIiIiKqqqru7u7u7u8zMzLu7u7u7u6qqqpmZmZmZmaqqqpmZmZmZmZmZmZmZmZmZmZmZmZmZmXd3d3d3d2ZmZnd3d3d3d3d3d3d3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVURERERERERERERERFVVVURERFVVVVVVVVVVVWZmZnd3d4iIiJmZmZmZmaqqqqqqqoiIiIiIiHd3d4iIiIiIiJmZmZmZmaqqqqqqqpmZmZmZmXd3d3d3d2ZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZlVVVWZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZnd3d4iIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d5mZmZmZmaqqqru7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqqqqqpmZmZmZmZmZmaqqqqqqqqqqqqqqqpmZmYiIiHd3d3d3d1VVVURERERERDMzMzMzMzMzMzMzM0RERERERERERERERFVVVWZmZmZmZnd3d2ZmZnd3d3d3d2ZmZnd3d3d3d2ZmZnd3d2ZmZmZmZlVVVWZmZlVVVVVVVVVVVURERERERERERDMzMzMzM0RERERERERERERERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVXd3d4iIiGZmZlVVVVVVVVVVVTMzMzMzMzMzM0RERDMzMzMzM0RERDMzM0RERDMzMzMzMzMzM0RERDMzM0RERERERERERERERFVVVWZmZlVVVURERERERERERDMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIiIiIiIiIjMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzM0RERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMyIiIhERERERESIiIiIiIiIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIjMzMyIiIjMzMzMzMyIiIiIiIhERESIiIjMzMyIiIiIiIiIiIiIiIiIiIhERESIiIiIiIhERESIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIjMzMzMzM0RERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIjMzM0RERERERFVVVWZmZnd3d2ZmZmZmZkRERERERERERERERERERERERERERFVVVWZmZnd3d4iIiIiIiIiIiGZmZlVVVVVVVVVVVVVVVYiIiMzMzP///+7u7v///+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7u7u7////u7u7////u7u7u7u7u7u7u7u7MzMy7u7vMzMy7u7u7u7uqqqqqqqq7u7vMzMzd3d3d3d3u7u7u7u7u7u7u7u7u7u7////////u7u7////u7u7u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3MzMzd3d3d3d3MzMzMzMzMzMzMzMzd3d3d3d3d3d3d3d3MzMzd3d3d3d3MzMy7u7uZmZl3d3d3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3dmZmZ3d3d3d3d3d3d3d3dmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZ3d3eIiIiZmZmZmZmZmZmqqqqZmZmqqqqqqqqqqqq7u7u7u7u7u7uqqqqZmZmZmZmIiIiIiIh3d3d3d3d3d3dmZmZmZmZmZmZmZmZVVVVmZmZmZmZEREREREREREQzMzMzMzNEREQzMzMzMzNERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3eZmZmqqqqqqqq7u7u7u7uqqqp3d3d3d3dmZmZVVVVVVVVVVVVEREQzMzNERERERERERERERERERERVVVVVVVVVVVVmZmZ3d3eZmZmqqqqqqqrMzMzd3d3MzMzd3d3MzMzMzMzMzMy7u7u7u7uqqqqZmZmqqqqZmZmqqqqZmZmIiIh3d3dmZmZmZmZVVVVVVVVVVVVVVVVERERERERERERERERERERERERERERVVVVEREREREQzMzNERERERERVVVVVVVVVVVVmZmZ3d3eIiIiZmZmqqqqZmZmZmZmIiIiIiIiIiIiIiIh3d3eIiIiZmZmqqqqqqqqZmZl3d3d3d3dmZmZVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVmZmZVVVVmZmZ3d3eIiIiZmZmIiIh3d3eIiIhmZmZ3d3d3d3eIiIiZmZmqqqqqqqqqqqqqqqqqqqq7u7u7u7u7u7u7u7u7u7uqqqqZmZmZmZmZmZmIiIiZmZmqqqqqqqqqqqqZmZmIiIiIiIh3d3dVVVVEREREREREREREREQzMzNEREQzMzNERERERERVVVVVVVVmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZVVVVmZmZ3d3d3d3dVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERVVVVERERVVVVVVVVmZmZ3d3dmZmZVVVVEREREREREREREREREREREREQzMzMzMzNEREREREREREREREREREREREREREQzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzMiIiIiIiIiIiIiIiIzMzMiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIzMzMzMzMiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIREREiIiIREREiIiIiIiIREREREREiIiIREREREREiIiIREREiIiIiIiIiIiIREREREREiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIREREiIiIREREREREREREiIiIREREiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIiIiIzMzMiIiIzMzMzMzMiIiIiIiIiIiIiIiIzMzMzMzNERERVVVVVVVVVVVVVVVVEREREREREREREREQzMzNERERVVVVmZmaIiIiZmZmZmZlmZmZVVVVERERERERERERERESZmZnd3d3u7u7////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u7u7u3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3du7u7qqqqmZmZmZmZiIiImZmZmZmZqqqqqqqqqqqqqqqqu7u7zMzMzMzMu7u7u7u7zMzM7u7u3d3dzMzMzMzM3d3dzMzM3d3dzMzM3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzM3d3dzMzMzMzMu7u7u7u7u7u7qqqqmZmZmZmZiIiId3d3d3d3d3d3ZmZmd3d3ZmZmd3d3ZmZmd3d3d3d3d3d3ZmZmd3d3d3d3d3d3iIiId3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmVVVVREREREREVVVVVVVVVVVVZmZmd3d3iIiIiIiImZmZqqqqu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7qqqqqqqqqqqqmZmZmZmZiIiIiIiIiIiId3d3ZmZmZmZmVVVVVVVVVVVVREREREREREREREREREREMzMzMzMzREREREREREREREREVVVVVVVVVVVVZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiImZmZqqqqu7u7u7u7qqqqiIiIiIiId3d3d3d3d3d3ZmZmREREREREREREREREREREVVVVREREVVVVVVVVVVVVZmZmd3d3d3d3iIiIqqqqu7u7u7u7zMzMzMzMzMzMzMzMzMzMu7u7qqqqmZmZiIiImZmZmZmZmZmZqqqqmZmZd3d3d3d3ZmZmVVVVREREREREREREREREREREREREMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzREREREREVVVVVVVVZmZmZmZmiIiIiIiIiIiIiIiImZmZmZmZiIiIiIiId3d3d3d3ZmZmd3d3iIiIiIiIiIiId3d3d3d3ZmZmVVVVVVVVREREREREREREREREREREREREVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmVVVVREREVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVd3d3iIiImZmZmZmZmZmZd3d3d3d3d3d3d3d3d3d3iIiImZmZmZmZqqqqqqqqqqqqu7u7qqqqu7u7u7u7qqqqqqqqmZmZmZmZmZmZiIiIiIiImZmZmZmZiIiImZmZiIiId3d3ZmZmVVVVVVVVREREMzMzREREMzMzMzMzREREREREREREREREZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmd3d3iIiId3d3ZmZmd3d3iIiIZmZmREREREREREREREREREREMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzREREVVVVVVVVVVVVREREVVVVREREREREMzMzIiIiMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzREREREREREREREREVVVVMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiERERIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERERERIiIiERERIiIiIiIiERERERERIiIiERERERERIiIiERERERERIiIiERERERERIiIiERERIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiERERERERIiIiIiIiERERIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERERERIiIiERERIiIiIiIiIiIiIiIiERERERERERERIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzREREREREREREMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREZmZmZmZmd3d3VVVVREREREREREREREREREREVVVVd3d3mZmZu7u77u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////+7u7u7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3czMzLu7u7u7u7u7u8zMzMzMzMzMzMzMzLu7u8zMzLu7u7u7u7u7u6qqqru7u8zMzMzMzMzMzMzMzMzMzMzMzN3d3d3d3czMzN3d3d3d3e7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3czMzMzMzMzMzLu7u6qqqqqqqqqqqpmZmYiIiIiIiJmZmZmZmZmZmZmZmZmZmZmZmYiIiHd3d3d3d3d3d3d3d3d3d2ZmZmZmZnd3d2ZmZnd3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVWZmZmZmZnd3d4iIiKqqqqqqqru7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqqqqqpmZmZmZmaqqqpmZmZmZmXd3d2ZmZmZmZkRERERERERERERERERERERERERERERERERERERERDMzM0RERERERERERGZmZmZmZnd3d3d3d4iIiIiIiJmZmZmZmYiIiIiIiIiIiHd3d4iIiIiIiJmZmaqqqqqqqpmZmZmZmZmZmZmZmXd3d1VVVWZmZlVVVVVVVURERFVVVVVVVURERFVVVVVVVWZmZmZmZmZmZnd3d4iIiIiIiKqqqqqqqru7u6qqqru7u6qqqqqqqpmZmYiIiIiIiIiIiIiIiJmZmYiIiIiIiIiIiHd3d3d3d2ZmZlVVVVVVVVVVVURERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERERERERERERERFVVVWZmZmZmZmZmZnd3d4iIiIiIiKqqqpmZmZmZmYiIiIiIiIiIiHd3d3d3d2ZmZmZmZmZmZmZmZnd3d3d3d1VVVVVVVURERDMzM0RERDMzM0RERERERFVVVURERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d2ZmZmZmZlVVVVVVVVVVVWZmZoiIiJmZmZmZmZmZmYiIiHd3d3d3d3d3d3d3d3d3d4iIiJmZmZmZmZmZmaqqqqqqqru7u7u7u7u7u6qqqqqqqpmZmZmZmYiIiIiIiIiIiIiIiJmZmZmZmZmZmYiIiHd3d2ZmZlVVVURERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVXd3d5mZmaqqqnd3d2ZmZmZmZnd3d2ZmZlVVVVVVVURERERERERERERERDMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzM0RERDMzMzMzMyIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzM0RERDMzMzMzMyIiIjMzMyIiIjMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIhERERERERERERERESIiIhERERERESIiIiIiIiIiIiIiIhERESIiIiIiIhERESIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERERERESIiIhERESIiIhERERERESIiIhERESIiIhERESIiIiIiIhERERERESIiIhERESIiIhERESIiIhERERERESIiIhERERERESIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIhERESIiIjMzMyIiIhERERERESIiIiIiIhERERERESIiIhERESIiIhERESIiIiIiIiIiIhERERERESIiIiIiIhERERERESIiIhERERERESIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMyIiIiIiIhERESIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIjMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMyIiIiIiIjMzMyIiIiIiIjMzMzMzMzMzM0RERERERERERERERERERERERDMzMzMzMzMzM0RERERERFVVVZmZmczMzO7u7v///////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7d3d3u7u7d3d3u7u7d3d3u7u7d3d3d3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7d3d3u7u7u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3MzMy7u7uqqqqqqqqqqqqZmZmZmZmZmZmIiIiIiIh3d3eIiIiIiIiZmZmZmZmZmZmZmZmqqqqqqqq7u7uqqqqZmZmIiIh3d3d3d3dmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZ3d3eIiIiZmZmqqqq7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7uqqqqqqqqqqqqqqqqqqqqqqqqqqqqZmZmIiIh3d3dmZmZVVVVVVVVERERERERERERERERERERERERERERERERERERmZmZmZmaIiIiIiIiIiIiZmZmZmZmZmZmZmZmZmZmIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZmZmZmqqqqZmZmIiIh3d3dmZmZ3d3dmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZ3d3eIiIiIiIiIiIiZmZmIiIiZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVEREREREREREQzMzNEREQzMzMzMzMzMzMzMzNERERERERERERERERERERVVVVVVVVmZmZmZmZ3d3eIiIiZmZmZmZmIiIiIiIiZmZmZmZmZmZmIiIhmZmZmZmZmZmZVVVVmZmZVVVVmZmZVVVVVVVVEREREREQzMzNERERERERVVVVERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVmZmZmZmZmZmZVVVVmZmZmZmZ3d3d3d3eIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3eIiIiIiIiIiIiZmZmZmZmqqqqqqqqqqqqqqqq7u7uqqqqqqqqZmZmZmZmZmZmZmZmZmZmIiIiZmZmZmZmZmZmZmZl3d3dmZmZEREREREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzNERERERERERERVVVVERERERERERERVVVVVVVV3d3eZmZl3d3dmZmZVVVVmZmZmZmZmZmZVVVVVVVVVVVVEREQzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIREREREREiIiIREREiIiIREREREREREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIREREiIiIREREREREiIiIREREiIiIREREREREREREiIiIREREREREREREiIiIiIiIiIiIzMzMiIiIzMzMiIiIREREiIiIREREREREREREiIiIREREREREiIiIREREREREREREREREiIiIREREREREREREiIiIiIiIiIiIREREiIiIREREREREREREiIiIREREiIiIREREiIiIREREiIiIREREREREiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIREREREREREREiIiIiIiIREREREREiIiIiIiIREREREREiIiIiIiIREREREREREREiIiIiIiIzMzMiIiIREREiIiIiIiIiIiIREREREREiIiIiIiIREREREREiIiIREREiIiIiIiIiIiIzMzMiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzNEREREREREREREREQzMzNERERERERVVVVVVVWIiIiqqqrd3d3////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////7u7u////////////////////////////////////7u7u////////////////7u7u////////////////////////7u7u////////////////7u7u////7u7u////7u7u////////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3d3d3dzMzMqqqqmZmZiIiIiIiIiIiIiIiId3d3d3d3iIiId3d3d3d3iIiImZmZiIiImZmZqqqqqqqqqqqqu7u7zMzMzMzMzMzMu7u7u7u7qqqqmZmZiIiId3d3d3d3VVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3iIiImZmZqqqqu7u7zMzMu7u7zMzMu7u7u7u7qqqqqqqqqqqqu7u7qqqqu7u7qqqqu7u7qqqqmZmZiIiId3d3d3d3ZmZmVVVVREREREREREREREREREREVVVVZmZmZmZmd3d3mZmZmZmZqqqqqqqqqqqqqqqqqqqqmZmZmZmZmZmZmZmZmZmZiIiIiIiIiIiId3d3iIiImZmZmZmZmZmZd3d3iIiImZmZiIiIiIiId3d3d3d3iIiIiIiId3d3ZmZmZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiIiIiIiIiImZmZiIiImZmZmZmZqqqqmZmZqqqqqqqqqqqqiIiId3d3d3d3ZmZmd3d3ZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREREREREREMzMzMzMzREREREREMzMzREREREREREREVVVVVVVVVVVVZmZmd3d3d3d3iIiIiIiImZmZmZmZqqqqqqqqqqqqiIiIiIiId3d3ZmZmVVVVVVVVREREREREVVVVVVVVREREREREREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3ZmZmVVVVVVVVZmZmZmZmd3d3iIiIiIiId3d3d3d3d3d3ZmZmd3d3d3d3iIiIiIiIiIiIiIiImZmZmZmZmZmZqqqqqqqqmZmZmZmZmZmZmZmZmZmZmZmZmZmZiIiIiIiImZmZqqqqqqqqmZmZVVVVREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREREREVVVVd3d3ZmZmVVVVZmZmVVVVZmZmZmZmVVVVREREMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERERERIiIiERERERERIiIiERERIiIiERERERERERERIiIiERERERERIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiMzMzMzMzIiIiIiIiMzMzIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiERERERERIiIiERERIiIiERERERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERERERIiIiIiIiERERERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERERERERERIiIiERERERERIiIiERERERERIiIiERERIiIiIiIiIiIiIiIiIiIiERERIiIiERERERERERERIiIiERERERERIiIiERERIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiERERERERERERERERIiIiERERIiIiIiIiIiIiERERIiIiERERERERIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzREREMzMzMzMzREREREREREREVVVVZmZmVVVVd3d3mZmZzMzM7u7u3d3d7u7u7u7u////////////////////////////////7u7u////////////////////////7u7u////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////+7u7v///////////+7u7v///////////////////////////////////////////////////////////////+7u7u7u7v///+7u7u7u7u7u7u7u7v///////+7u7v///+7u7v///+7u7v///+7u7v///+7u7v///+7u7v///+7u7v///+7u7v///+7u7u7u7v///+7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzN3d3czMzMzMzN3d3d3d3d3d3d3d3d3d3e7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3czMzKqqqoiIiHd3d3d3d2ZmZnd3d3d3d3d3d3d3d2ZmZnd3d4iIiIiIiJmZmZmZmaqqqqqqqqqqqru7u8zMzLu7u8zMzLu7u8zMzLu7u8zMzLu7u6qqqpmZmaqqqoiIiIiIiGZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiJmZmZmZmaqqqru7u7u7u7u7u7u7u6qqqqqqqqqqqqqqqqqqqoiIiJmZmaqqqqqqqqqqqpmZmZmZmYiIiHd3d2ZmZlVVVVVVVVVVVVVVVVVVVWZmZnd3d4iIiJmZmaqqqru7u7u7u6qqqpmZmZmZmaqqqqqqqqqqqpmZmZmZmZmZmZmZmYiIiIiIiHd3d3d3d3d3d2ZmZmZmZnd3d4iIiJmZmZmZmYiIiIiIiJmZmaqqqpmZmZmZmXd3d2ZmZnd3d2ZmZnd3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiJmZmYiIiJmZmaqqqqqqqqqqqqqqqpmZmXd3d3d3d2ZmZnd3d3d3d3d3d2ZmZmZmZnd3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVURERERERERERERERERERERERFVVVVVVVVVVVVVVVWZmZlVVVWZmZnd3d3d3d4iIiIiIiJmZmaqqqqqqqqqqqpmZmaqqqpmZmZmZmXd3d2ZmZmZmZlVVVURERERERERERERERERERERERFVVVURERERERERERERERERERERERERERFVVVURERFVVVVVVVURERGZmZlVVVWZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZnd3d3d3d3d3d3d3d2ZmZnd3d2ZmZnd3d3d3d4iIiHd3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiJmZmZmZmZmZmZmZmZmZmZmZmYiIiHd3d6qqqru7u6qqqnd3d2ZmZmZmZlVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzM0RERFVVVURERERERERERERERERERDMzMyIiIiIiIiIiIhERESIiIhERESIiIhERERERERERERERERERERERERERERERESIiIhERERERERERESIiIhERESIiIhERESIiIhERERERESIiIhERESIiIhERESIiIhERERERESIiIhERESIiIjMzMzMzMyIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIjMzMzMzMyIiIiIiIjMzMyIiIiIiIhERESIiIhERESIiIhERERERESIiIhERESIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIhERESIiIhERERERERERESIiIhERERERESIiIhERESIiIiIiIiIiIiIiIhERERERERERESIiIhERESIiIhERERERESIiIhERERERESIiIhERERERERERESIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIhERERERESIiIhERESIiIiIiIhERERERESIiIiIiIiIiIiIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERDMzM0RERERERERERERERFVVVVVVVVVVVWZmZmZmZoiIiJmZmZmZmaqqqszMzN3d3e7u7u7u7u7u7v///////////////////////////////+7u7v///////////////////+7u7v///////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////u7u7u7u7d3d3u7u7u7u7////d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7////u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3MzMzd3d3MzMzd3d3MzMzMzMzd3d3MzMzMzMzd3d3d3d3d3d3u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3MzMy7u7uZmZl3d3d3d3dmZmZ3d3d3d3d3d3d3d3dmZmZ3d3d3d3eZmZmqqqqZmZmZmZmqqqq7u7u7u7u7u7vMzMzMzMzMzMy7u7vMzMy7u7u7u7uqqqqqqqqqqqq7u7uqqqqZmZmZmZmIiIh3d3dmZmZmZmZERERVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZ3d3d3d3eIiIiIiIiZmZmZmZmqqqqqqqqZmZmZmZmZmZmZmZmIiIiZmZmIiIiZmZmZmZmqqqqqqqq7u7uqqqqqqqqqqqqZmZmZmZmZmZmZmZmZmZmZmZmZmZmqqqqqqqqZmZmZmZmIiIh3d3d3d3dmZmZmZmZmZmZ3d3d3d3eIiIiZmZmqqqqqqqqZmZmqqqqZmZmZmZmZmZmZmZmZmZmZmZmZmZmIiIh3d3d3d3d3d3d3d3dmZmZVVVVVVVVmZmZ3d3d3d3eIiIiIiIiIiIiIiIiZmZmZmZmZmZmIiIiIiIiIiIiIiIhmZmZmZmZmZmZ3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZmqqqqqqqqZmZmIiIiIiIh3d3d3d3dmZmZ3d3dmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3dVVVVmZmZVVVVVVVVVVVVERERERERVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZ3d3d3d3eIiIiIiIiIiIiZmZmZmZmZmZmZmZmqqqqqqqqqqqqZmZmZmZmZmZl3d3dmZmZVVVVEREREREQzMzNERERERERERERERERERERERERERERERERERERERERVVVVERERERERVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZVVVVERERVVVVmZmZmZmZmZmZ3d3dmZmZmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZ3d3dmZmZ3d3d3d3eIiIh3d3eIiIh3d3eIiIiIiIh3d3d3d3d3d3d3d3eIiIiIiIiIiIh3d3dmZmZVVVVEREREREQzMzMzMzNEREQzMzMzMzNEREQzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMiIiIiIiIiIiIiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIREREREREREREREREiIiIREREiIiIREREiIiIREREREREiIiIREREREREiIiIiIiIiIiIiIiIREREiIiIREREiIiIiIiIzMzMiIiIzMzMzMzMiIiIiIiIiIiIzMzMiIiIiIiIzMzMiIiIzMzMzMzMiIiIzMzMzMzMiIiIiIiIiIiIiIiIREREREREiIiIREREiIiIREREREREiIiIREREREREREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIiIiIREREREREiIiIREREiIiIREREREREiIiIREREiIiIREREREREiIiIREREiIiIREREREREiIiIREREiIiIREREiIiIREREREREREREREREiIiIREREREREiIiIiIiIiIiIiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIREREREREiIiIREREiIiIREREREREiIiIiIiIREREREREiIiIREREREREiIiIiIiIREREREREiIiIREREREREzMzMzMzMiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMzMzMzMzNERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmaIiIiIiIiZmZmqqqq7u7vMzMzd3d3u7u7u7u7u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////7u7u7u7u////7u7u////7u7u3d3d3d3du7u7zMzMzMzMzMzMqqqqqqqqu7u7u7u7zMzM3d3dzMzMzMzMzMzM3d3d3d3d3d3d7u7u7u7u3d3d7u7u3d3d7u7u7u7u3d3d7u7u7u7u////7u7u7u7u////7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u7u7u3d3d7u7u7u7u3d3d7u7u3d3dzMzMu7u7iIiId3d3d3d3ZmZmd3d3ZmZmd3d3d3d3iIiIiIiIiIiImZmZqqqqmZmZqqqqqqqqu7u7mZmZqqqqu7u7u7u7zMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7qqqqqqqqqqqqqqqqmZmZqqqqmZmZmZmZiIiId3d3ZmZmVVVVVVVVREREVVVVREREVVVVREREZmZmZmZmZmZmZmZmd3d3iIiImZmZqqqqqqqqu7u7u7u7u7u7qqqqqqqqmZmZqqqqmZmZmZmZmZmZiIiImZmZmZmZqqqqqqqqqqqqqqqqmZmZmZmZmZmZiIiIiIiIiIiImZmZmZmZqqqqqqqqqqqqmZmZmZmZiIiIiIiIiIiId3d3d3d3d3d3iIiId3d3iIiIiIiImZmZiIiImZmZmZmZmZmZmZmZmZmZmZmZiIiId3d3d3d3d3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3ZmZmd3d3iIiIiIiIiIiIiIiImZmZmZmZmZmZiIiId3d3d3d3ZmZmZmZmZmZmd3d3iIiId3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiImZmZmZmZiIiImZmZiIiId3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3ZmZmZmZmVVVVVVVVZmZmVVVVVVVVVVVVZmZmd3d3d3d3d3d3d3d3iIiIiIiIiIiImZmZmZmZmZmZmZmZiIiImZmZmZmZmZmZqqqqmZmZmZmZmZmZmZmZd3d3ZmZmVVVVREREREREMzMzREREREREREREMzMzREREREREVVVVREREREREREREREREREREREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmVVVVZmZmd3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3ZmZmZmZmZmZmd3d3ZmZmVVVVVVVVREREREREMzMzREREMzMzREREMzMzREREMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiIiIiERERERERIiIiERERERERIiIiERERIiIiERERIiIiERERERERIiIiERERERERERERIiIiERERERERERERERERIiIiERERIiIiERERERERERERIiIiERERERERIiIiERERERERIiIiERERERERERERIiIiIiIiIiIiERERIiIiIiIiMzMzIiIiIiIiMzMzREREMzMzIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERERERIiIiIiIiERERERERIiIiERERIiIiERERIiIiERERIiIiERERERERIiIiERERIiIiERERERERERERIiIiERERERERIiIiERERERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERERERERERIiIiERERERERIiIiERERIiIiIiIiIiIiERERIiIiERERIiIiERERERERIiIiIiIiERERIiIiIiIiMzMzIiIiIiIiERERIiIiERERIiIiERERIiIiERERERERIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiERERERERIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERERERERERIiIiERERIiIiIiIiMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiERERERERERERERERIiIiMzMzIiIiERERIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzREREMzMzREREREREREREVVVVREREREREVVVVVVVVZmZmZmZmd3d3iIiImZmZqqqqzMzM3d3d3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////+7u7u7u7u7u7t3d3e7u7u7u7u7u7t3d3d3d3d3d3czMzMzMzMzMzLu7u8zMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3d3d3e7u7t3d3e7u7t3d3d3d3d3d3e7u7u7u7u7u7u7u7v///+7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3czMzMzMzMzMzMzMzMzMzMzMzN3d3czMzN3d3e7u7t3d3d3d3czMzN3d3d3d3d3d3czMzMzMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u7u7u8zMzLu7u5mZmXd3d3d3d3d3d2ZmZmZmZmZmZoiIiIiIiIiIiJmZmaqqqqqqqqqqqqqqqqqqqru7u6qqqqqqqqqqqru7u7u7u7u7u8zMzMzMzLu7u6qqqru7u6qqqru7u6qqqqqqqqqqqpmZmZmZmYiIiJmZmZmZmZmZmZmZmYiIiHd3d4iIiHd3d2ZmZlVVVVVVVURERERERFVVVVVVVWZmZnd3d3d3d4iIiKqqqru7u6qqqqqqqqqqqru7u6qqqqqqqqqqqqqqqru7u6qqqqqqqpmZmYiIiIiIiIiIiIiIiJmZmZmZmZmZmZmZmYiIiHd3d3d3d3d3d3d3d4iIiJmZmZmZmZmZmZmZmaqqqqqqqpmZmaqqqpmZmZmZmZmZmYiIiIiIiHd3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d2ZmZlVVVVVVVURERFVVVURERERERFVVVURERFVVVWZmZlVVVWZmZnd3d3d3d2ZmZnd3d5mZmZmZmZmZmZmZmYiIiIiIiHd3d2ZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d4iIiIiIiHd3d2ZmZmZmZmZmZnd3d4iIiIiIiHd3d2ZmZnd3d1VVVWZmZlVVVWZmZmZmZmZmZnd3d4iIiJmZmZmZmZmZmZmZmaqqqqqqqpmZmZmZmZmZmYiIiIiIiIiIiJmZmZmZmZmZmZmZmZmZmZmZmXd3d2ZmZmZmZkRERERERDMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERERERFVVVURERFVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZmZmZoiIiHd3d2ZmZmZmZmZmZlVVVVVVVVVVVURERERERDMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMyIiIiIiIiIiIhERESIiIjMzMyIiIhERESIiIiIiIhERERERESIiIhERERERESIiIhERERERERERESIiIhERERERESIiIhERESIiIhERESIiIhERERERESIiIhERESIiIhERERERERERESIiIhERESIiIhERESIiIhERERERERERESIiIhERERERESIiIhERESIiIiIiIiIiIiIiIhERESIiIiIiIiIiIhERESIiIjMzMyIiIjMzMyIiIjMzMzMzMyIiIiIiIiIiIhERERERERERERERERERESIiIiIiIhERESIiIiIiIhERESIiIiIiIiIiIhERESIiIhERESIiIhERESIiIhERERERESIiIhERERERESIiIhERERERESIiIhERESIiIhERESIiIhERERERESIiIhERERERESIiIhERESIiIhERERERESIiIiIiIiIiIhERERERESIiIhERESIiIhERESIiIhERERERESIiIhERESIiIiIiIiIiIhERESIiIhERERERESIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIhERERERESIiIhERESIiIhERERERESIiIhERERERESIiIhERESIiIhERERERESIiIhERERERESIiIhERESIiIhERESIiIhERERERESIiIiIiIhERERERESIiIhERERERESIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIhERESIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIhERERERERERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMyIiIjMzMzMzM0RERERERFVVVURERERERERERERERFVVVWZmZmZmZmZmZnd3d3d3d5mZmaqqqqqqqszMzMzMzO7u7u7u7v///+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////u7u7////u7u7u7u7////u7u7////u7u7////u7u7u7u7d3d3u7u7d3d3u7u7u7u7u7u7////u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7d3d3d3d3d3d3u7u7d3d3u7u7u7u7d3d3u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3d3d3MzMzMzMzMzMzd3d3MzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7uqqqqqqqqZmZmZmZmZmZmZmZmIiIiZmZmZmZmIiIh3d3d3d3dmZmZmZmZmZmZmZmZ3d3eIiIiZmZmIiIiZmZmqqqq7u7uqqqq7u7u7u7u7u7u7u7u7u7u7u7u7u7uqqqq7u7u7u7u7u7uqqqrMzMy7u7u7u7uqqqqqqqqZmZmZmZmZmZmIiIiIiIiIiIiIiIiIiIiIiIiZmZmZmZmqqqqqqqqZmZmIiIiIiIhmZmZVVVVVVVVVVVVVVVVmZmZ3d3eIiIiZmZmqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqq7u7uqqqqqqqqqqqqqqqqZmZmIiIiIiIh3d3eIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3eIiIhmZmZ3d3d3d3eIiIiZmZmZmZmqqqq7u7u7u7u7u7uqqqqqqqqZmZmIiIh3d3d3d3eIiIiIiIiIiIiIiIh3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVERERERERVVVVERERERERVVVVVVVVmZmZVVVVmZmaIiIiIiIiZmZmZmZmZmZmIiIiIiIh3d3eIiIh3d3dmZmZVVVVVVVVmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIh3d3eIiIh3d3dmZmZVVVVmZmZmZmZmZmZ3d3eIiIiIiIh3d3d3d3dmZmZ3d3dmZmZ3d3d3d3d3d3d3d3eZmZmZmZmZmZmqqqqqqqqqqqq7u7uqqqqZmZmIiIiIiIiZmZmIiIiZmZmZmZmqqqqZmZmZmZmIiIh3d3dmZmZmZmZEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZmZmZVVVVVVVVVVVVVVVVERERERERERERERERVVVVVVVVEREREREQzMzNERERERERVVVVVVVVmZmZmZmZVVVVVVVVVVVVERERVVVVEREQzMzNEREQzMzMzMzMzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIREREiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIREREREREiIiIREREREREiIiIREREREREiIiIREREiIiIREREiIiIREREiIiIREREREREiIiIREREREREREREiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIiIiIzMzMiIiIREREiIiIiIiIiIiIREREREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIREREiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIREREREREREREREREREREiIiIREREREREiIiIREREREREiIiIREREREREiIiIREREiIiIREREiIiIiIiIREREREREREREiIiIREREREREiIiIREREiIiIREREiIiIREREiIiIREREREREREREiIiIREREiIiIiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIREREREREREREiIiIREREiIiIiIiIREREREREiIiIiIiIREREiIiIiIiIiIiIREREREREiIiIREREREREiIiIREREREREiIiIREREREREREREiIiIREREREREiIiIREREiIiIiIiIiIiIREREREREiIiIREREREREREREiIiIREREiIiIREREiIiIREREREREiIiIiIiIiIiIiIiIzMzMREREiIiIREREREREREREiIiIREREiIiIREREREREREREiIiIREREiIiIiIiIiIiIREREREREREREiIiIREREREREiIiIREREREREiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMiIiIiIiIzMzMiIiIzMzMzMzNVVVVVVVVERERERERVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZ3d3eIiIiIiIiZmZmqqqrMzMzMzMzd3d3u7u7u7u7////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3d3d3d7u7u7u7u7u7u7u7u////////////////////7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d7u7u7u7u3d3d7u7u3d3d7u7u7u7u7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d7u7u3d3d3d3d3d3dzMzMzMzMu7u7zMzMzMzMzMzMzMzM3d3dzMzMzMzM3d3d3d3d3d3dzMzMzMzMu7u7qqqqqqqqqqqqqqqqqqqqmZmZmZmZmZmZqqqqiIiIiIiId3d3iIiId3d3d3d3ZmZmZmZmZmZmZmZmd3d3mZmZmZmZmZmZmZmZqqqqzMzMu7u7u7u7u7u7u7u7zMzMu7u7u7u7u7u7u7u7zMzMzMzMu7u7u7u7u7u7u7u7u7u7zMzMu7u7u7u7qqqqiIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiImZmZmZmZqqqqqqqqqqqqqqqqmZmZiIiId3d3d3d3ZmZmd3d3iIiImZmZmZmZmZmZmZmZmZmZmZmZqqqqmZmZqqqqqqqqqqqqqqqqu7u7qqqqqqqqmZmZqqqqmZmZiIiIiIiId3d3d3d3d3d3d3d3ZmZmZmZmd3d3d3d3iIiIZmZmZmZmVVVVd3d3ZmZmd3d3iIiImZmZqqqqqqqqu7u7u7u7u7u7mZmZmZmZiIiIiIiId3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiImZmZd3d3ZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3iIiIiIiIiIiId3d3ZmZmZmZmZmZmZmZmZmZmd3d3d3d3iIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmd3d3d3d3iIiImZmZmZmZmZmZmZmZqqqqqqqqqqqqqqqqmZmZmZmZiIiIiIiIiIiIiIiIiIiImZmZmZmZmZmZiIiId3d3ZmZmVVVVVVVVREREREREREREMzMzMzMzMzMzMzMzREREMzMzMzMzREREREREVVVVVVVVVVVVZmZmVVVVZmZmVVVVZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREVVVVREREMzMzREREMzMzREREREREREREREREREREREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzIiIiIiIiERERERERERERIiIiERERIiIiIiIiIiIiERERERERERERIiIiERERERERERERERERIiIiERERIiIiERERERERIiIiERERERERIiIiERERERERIiIiERERIiIiERERERERERERIiIiERERERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERERERIiIiERERERERIiIiIiIiIiIiIiIiERERERERERERERERERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiERERERERIiIiERERERERIiIiERERERERIiIiIiIiERERIiIiERERIiIiIiIiERERIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiERERIiIiIiIiERERIiIiIiIiERERIiIiERERERERERERERERIiIiERERIiIiERERERERERERIiIiERERERERERERERERIiIiIiIiIiIiERERIiIiERERIiIiIiIiERERERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiERERERERIiIiERERIiIiERERERERERERIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiIiIiERERIiIiERERIiIiEREREREA//8AABEiIiIiIiIiIiIiIiIiIiIREREiIiIREREREREiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzNVVVVVVVVEREQzMzNERERERERERERERERERERVVVVVVVVVVVVmZmZmZmZ3d3d3d3eIiIiZmZmqqqq7u7vMzMzd3d3d3d3u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3dzMzMzMzMzMzMzMzM3d3d3d3d7u7u7u7u7u7u7u7u////7u7u7u7u////7u7u7u7u////7u7u7u7u7u7u7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u////7u7u7u7u7u7u3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMu7u7qqqqqqqqqqqqmZmZmZmZmZmZqqqqmZmZmZmZmZmZmZmZmZmZiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmiIiIiIiIiIiImZmZqqqqu7u7zMzMu7u7zMzMzMzMzMzMu7u7u7u7zMzMzMzMzMzMzMzMu7u7zMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7mZmZmZmZiIiId3d3d3d3VVVVVVVVZmZmZmZmZmZmd3d3d3d3iIiIiIiIiIiIqqqqqqqqu7u7u7u7u7u7u7u7u7u7mZmZmZmZiIiImZmZmZmZmZmZmZmZmZmZqqqqqqqqmZmZqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqmZmZiIiImZmZiIiIiIiIZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmVVVVZmZmd3d3iIiIiIiIiIiIqqqqqqqqu7u7u7u7qqqqqqqqiIiId3d3d3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiImZmZqqqqmZmZiIiIiIiIiIiIiIiId3d3d3d3ZmZmVVVVZmZmVVVVZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmd3d3ZmZmd3d3d3d3d3d3ZmZmVVVVZmZmVVVVZmZmZmZmZmZmd3d3iIiIiIiIiIiId3d3d3d3iIiIiIiIiIiIiIiImZmZmZmZmZmZmZmZqqqqqqqqqqqqmZmZmZmZiIiIiIiId3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiIZmZmZmZmVVVVVVVVVVVVMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREMzMzREREREREVVVVREREREREVVVVVVVVVVVVVVVVVVVVZmZmd3d3iIiId3d3d3d3ZmZmVVVVVVVVZmZmd3d3d3d3ZmZmZmZmVVVVREREREREREREREREREREMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiERERIiIiERERIiIiERERERERIiIiIiIiIiIiIiIiERERERERERERIiIiERERIiIiERERIiIiERERERERIiIiERERERERIiIiERERERERIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiERERERERERERERERIiIiERERERERERERIiIiERERIiIiERERERERIiIiIiIiERERIiIiMzMzMzMzIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiERERERERIiIiMzMzIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiERERERERIiIiIiIiIiIiIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiERERERERIiIiERERERERERERERERIiIiERERERERERERIiIiERERERERIiIiERERIiIiERERERERIiIiIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERERERIiIiERERERERERERIiIiERERIiIiIiIiIiIiERERERERERERIiIiERERERERIiIiERERIiIiERERIiIiERERERERIiIiERERIiIiMzMzIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERERERIiIiERERERERIiIiERERERERIiIiIiIiIiIiERERERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzMzMzREREMzMzMzMzMzMzMzMzREREMzMzREREREREVVVVREREVVVVVVVVVVVVZmZmZmZmd3d3d3d3iIiIiIiIqqqqzMzM3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////+7u7v///////////////////////////+7u7v///+7u7v///+7u7u7u7t3d3d3d3d3d3czMzMzMzN3d3czMzMzMzMzMzN3d3czMzN3d3d3d3e7u7u7u7u7u7v///+7u7u7u7v///+7u7u7u7u7u7u7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7v///+7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7u7u7t3d3e7u7t3d3e7u7u7u7u7u7u7u7t3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3czMzKqqqpmZmYiIiIiIiHd3d4iIiJmZmZmZmZmZmYiIiJmZmYiIiHd3d4iIiIiIiJmZmZmZmYiIiIiIiIiIiJmZmYiIiIiIiIiIiHd3d5mZmZmZmaqqqqqqqru7u6qqqru7u7u7u7u7u6qqqru7u7u7u7u7u7u7u7u7u6qqqru7u6qqqqqqqqqqqqqqqpmZmZmZmZmZmYiIiHd3d3d3d3d3d2ZmZlVVVWZmZlVVVVVVVWZmZmZmZlVVVWZmZmZmZoiIiIiIiIiIiKqqqru7u7u7u7u7u8zMzMzMzLu7u6qqqru7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqru7u7u7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqpmZmZmZmZmZmYiIiHd3d1VVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d4iIiKqqqru7u7u7u7u7u6qqqqqqqoiIiHd3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVURERERERERERFVVVVVVVVVVVURERFVVVVVVVVVVVVVVVWZmZnd3d2ZmZnd3d3d3d4iIiIiIiKqqqqqqqpmZmaqqqqqqqqqqqqqqqqqqqpmZmYiIiHd3d2ZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZlVVVWZmZmZmZlVVVWZmZmZmZnd3d2ZmZmZmZnd3d2ZmZmZmZlVVVVVVVWZmZmZmZnd3d4iIiIiIiIiIiIiIiHd3d4iIiIiIiJmZmYiIiJmZmYiIiJmZmYiIiJmZmZmZmZmZmZmZmYiIiJmZmYiIiIiIiIiIiIiIiHd3d4iIiHd3d3d3d3d3d2ZmZmZmZlVVVURERERERDMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERERERERERERERERERERERERERERERERERFVVVVVVVXd3d3d3d2ZmZnd3d3d3d3d3d1VVVWZmZnd3d3d3d2ZmZmZmZmZmZlVVVURERDMzM0RERDMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIhERESIiIhERERERESIiIhERESIiIjMzMyIiIhERESIiIhERESIiIhERESIiIhERESIiIhERERERESIiIhERERERESIiIhERERERESIiIhERESIiIhERESIiIhERESIiIhERERERERERERERESIiIhERESIiIhERESIiIhERESIiIhERESIiIhERERERESIiIiIiIhERERERESIiIiIiIhERETMzMyIiIiIiIiIiIhERESIiIiIiIhERESIiIhERESIiIhERESIiIiIiIhERESIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMyIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIhERERERESIiIhERESIiIiIiIhERERERERERESIiIiIiIjMzMyIiIiIiIhERERERESIiIhERERERERERESIiIhERESIiIhERESIiIhERERERESIiIhERERERESIiIhERERERESIiIhERESIiIiIiIhERERERERERESIiIhERERERERERERERESIiIiIiIiIiIhERESIiIhERERERERERESIiIiIiIhERERERERERESIiIiIiIhERERERESIiIiIiIhERESIiIhERERERERERESIiIhERESIiIhERESIiIhERERERESIiIhERERERERERERERERERESIiIhERERERESIiIiIiIiIiIhERESIiIhERESIiIhERERERESIiIhERERERESIiIhERESIiIhERERERESIiIhERESIiIhERERERESIiIiIiIiIiIhERESIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERETMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERFVVVVVVVWZmZlVVVWZmZmZmZnd3d4iIiIiIiKqqqszMzMzMzO7u7u7u7u7u7v///+7u7v///////////////+7u7v///////////////+7u7v///////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////u7u7////////u7u7////////////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3u7u7d3d3d3d3MzMzMzMzMzMzd3d3d3d3d3d3d3d3u7u7u7u7u7u7////////u7u7u7u7u7u7////u7u7////u7u7////u7u7////u7u7u7u7u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3MzMzd3d3d3d3d3d3MzMzd3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d27u7uZmZl3d3eIiIiIiIh3d3eIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3eIiIiZmZmIiIiZmZmIiIiZmZmZmZmZmZmZmZmIiIiZmZmZmZmqqqqZmZmqqqqZmZmqqqqqqqq7u7uqqqqqqqq7u7uqqqqqqqqqqqqqqqqqqqqqqqqZmZmIiIiIiIh3d3d3d3dmZmZ3d3d3d3dmZmZmZmZmZmZVVVVmZmZVVVVmZmZVVVVVVVVmZmZmZmZmZmZ3d3eIiIiIiIiZmZmqqqqqqqq7u7u7u7u7u7u7u7vMzMy7u7u7u7u7u7uqqqqqqqqqqqqZmZmqqqqqqqqZmZmqqqqqqqqZmZmZmZmqqqqZmZmqqqqZmZmZmZmIiIh3d3dmZmZVVVVVVVVVVVVmZmZVVVVVVVVVVVVERERVVVVmZmZmZmZ3d3d3d3dmZmZ3d3d3d3eIiIiZmZmZmZmqqqq7u7u7u7uqqqqZmZmIiIh3d3dmZmZVVVVVVVVERERVVVVERERVVVVERERERERERERERERERERERERERERERERVVVVERERVVVVVVVVmZmZmZmZ3d3d3d3d3d3eZmZmqqqqqqqq7u7uqqqq7u7u7u7uqqqq7u7u7u7uZmZmIiIh3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZ3d3d3d3dmZmZmZmZVVVVVVVVVVVVmZmZmZmZ3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIiZmZmZmZmZmZmIiIiIiIiIiIiIiIiIiIiZmZmIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZVVVVVVVVEREREREQzMzMzMzNEREREREREREREREREREREREREREREREQzMzNEREREREQzMzNERERERERERERVVVVERERVVVV3d3eIiIh3d3dmZmZVVVVmZmZVVVVEREREREREREQzMzMzMzMiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIREREREREREREiIiIREREiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREREREREREREREiIiIREREiIiIREREiIiIREREREREiIiIREREREREiIiIREREREREiIiIiIiIREREiIiIiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIREREREREiIiIREREiIiIREREREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIREREREREiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIREREREREREREREREiIiIREREiIiIREREREREiIiIiIiIiIiIREREiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIiIiIREREREREREREREREiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIREREiIiIREREREREiIiIREREREREiIiIiIiIREREiIiIREREREREiIiIREREREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIiIiIREREREREREREiIiIREREREREiIiIREREiIiIREREiIiIREREiIiIREREiIiIREREiIiIiIiIzMzMREREiIiIREREiIiIREREiIiIiIiIREREREREREREREREiIiIREREiIiIREREiIiIREREiIiIREREiIiIzMzMiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIREREzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzNEREQzMzNERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZ3d3eIiIiZmZm7u7vMzMzd3d3u7u7////////u7u7////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3dzMzM3d3dzMzM3d3d3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3dzMzMzMzMzMzMzMzM3d3d3d3d3d3d3d3d7u7u3d3d7u7u3d3d7u7u7u7u7u7u7u7u////////7u7u////////7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3dzMzMu7u7u7u7u7u7u7u7u7u7zMzMzMzM3d3d3d3d3d3d7u7u3d3d3d3d7u7u3d3d3d3d3d3dzMzMqqqqmZmZmZmZiIiIiIiIiIiId3d3iIiIiIiId3d3d3d3ZmZmd3d3ZmZmZmZmZmZmd3d3d3d3ZmZmd3d3d3d3iIiImZmZqqqqmZmZmZmZqqqqqqqqmZmZqqqqmZmZmZmZmZmZqqqqmZmZmZmZmZmZqqqqqqqqu7u7u7u7zMzMu7u7qqqqmZmZiIiId3d3d3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3iIiImZmZmZmZqqqqqqqqu7u7u7u7u7u7zMzMzMzMzMzMu7u7u7u7qqqqmZmZmZmZmZmZmZmZiIiIiIiImZmZmZmZmZmZmZmZmZmZiIiId3d3ZmZmVVVVVVVVREREREREREREREREREREREREVVVVVVVVVVVVZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiImZmZmZmZmZmZmZmZmZmZiIiId3d3d3d3VVVVVVVVVVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmd3d3d3d3mZmZmZmZu7u7u7u7zMzMzMzMzMzMzMzMzMzMu7u7u7u7qqqqmZmZd3d3d3d3VVVVVVVVVVVVREREVVVVREREREREVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmd3d3d3d3iIiIiIiIiIiIiIiImZmZmZmZiIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3iIiId3d3d3d3d3d3ZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmVVVVREREVVVVMzMzMzMzREREREREREREREREREREREREMzMzREREMzMzMzMzMzMzMzMzREREMzMzREREMzMzREREVVVVd3d3VVVVVVVVVVVVREREREREIiIiIiIiMzMzIiIiIiIiERERERERIiIiIiIiIiIiERERIiIiIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiMzMzIiIiIiIiERERERERIiIiERERMzMzIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiERERERERIiIiERERIiIiIiIiIiIiERERERERIiIiERERIiIiERERIiIiERERERERERERERERIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiERERERERERERIiIiERERERERIiIiERERIiIiERERERERIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiERERIiIiIiIiMzMzIiIiMzMzIiIiMzMzERERERERIiIiERERERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiERERIiIiERERIiIiERERERERERERIiIiERERERERERERIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiERERERERIiIiIiIiERERIiIiERERIiIiERERERERERERERERERERERERIiIiERERERERIiIiERERERERIiIiIiIiERERIiIiERERERERERERIiIiERERERERIiIiERERERERIiIiERERERERERERERERERERIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERERERIiIiERERIiIiIiIiIiIiIiIiERERIiIiIiIiERERERERIiIiERERERERIiIiERERERERIiIiERERERERIiIiIiIiIiIiIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiIiIiERERIiIiERERIiIiERERERERERERIiIiIiIiIiIiIiIiERERERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzMzMzMzMzVVVVREREREREREREREREVVVVVVVVVVVVZmZmd3d3d3d3mZmZmZmZqqqqzMzM7u7u7u7u////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////+7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3czMzN3d3czMzMzMzMzMzN3d3d3d3d3d3d3d3e7u7u7u7u7u7u7u7t3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7u7u7u7u7u7u7v///////////////+7u7v///+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzLu7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqru7u8zMzMzMzMzMzN3d3d3d3czMzN3d3czMzMzMzMzMzKqqqpmZmZmZmYiIiIiIiIiIiIiIiJmZmYiIiIiIiHd3d3d3d3d3d1VVVVVVVWZmZmZmZlVVVVVVVVVVVWZmZnd3d3d3d4iIiIiIiJmZmZmZmZmZmZmZmaqqqru7u6qqqqqqqru7u6qqqqqqqoiIiJmZmaqqqqqqqru7u7u7u6qqqqqqqoiIiIiIiHd3d2ZmZmZmZlVVVVVVVVVVVVVVVURERERERERERERERERERFVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d4iIiIiIiJmZmZmZmaqqqqqqqqqqqszMzMzMzMzMzMzMzMzMzLu7u6qqqpmZmZmZmYiIiIiIiIiIiIiIiIiIiIiIiHd3d2ZmZlVVVVVVVURERERERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d2ZmZlVVVVVVVWZmZmZmZnd3d4iIiIiIiIiIiJmZmZmZmZmZmYiIiGZmZmZmZlVVVURERERERERERFVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZnd3d3d3d3d3d4iIiJmZmaqqqru7u7u7u93d3czMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u5mZmYiIiHd3d1VVVVVVVURERERERDMzM0RERERERERERERERERERFVVVVVVVVVVVWZmZlVVVVVVVURERFVVVVVVVVVVVWZmZmZmZnd3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZnd3d2ZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERERERDMzM0RERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIhERESIiIhERESIiIhERESIiIhERERERESIiIhERESIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIhERERERESIiIiIiIiIiIiIiIhERESIiIhERERERERERESIiIhERESIiIhERERERERERESIiIhERERERESIiIhERERERESIiIhERERERERERESIiIhERESIiIhERESIiIhERERERESIiIhERERERESIiIhERERERESIiIhERESIiIhERERERESIiIhERESIiIhERERERESIiIhERERERERERESIiIhERESIiIhERESIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIhERERERESIiIhERERERESIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIhERESIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERERERESIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIhERESIiIiIiIiIiIhERESIiIhERERERERERESIiIhERERERESIiIhERERERESIiIiIiIhERESIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIhERERERESIiIhERERERESIiIiIiIiIiIhERESIiIhERERERESIiIiIiIhERESIiIhERERERERERERERERERERERESIiIhERESIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzM0RERERERERERDMzMzMzM0RERFVVVVVVVVVVVVVVVWZmZnd3d3d3d5mZmaqqqru7u8zMzN3d3e7u7u7u7v///////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7////////////u7u7////////////u7u7////////////u7u7////u7u7u7u7d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3MzMzd3d3d3d3d3d3u7u7d3d3u7u7d3d3u7u7u7u7d3d3d3d3MzMzd3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7////u7u7u7u7d3d3u7u7u7u7u7u7d3d3d3d3MzMzMzMzMzMzMzMy7u7u7u7u7u7uqqqqqqqq7u7uqqqqqqqqZmZmqqqqqqqqqqqq7u7u7u7u7u7uqqqq7u7uqqqqZmZmqqqqZmZmZmZmZmZmIiIiIiIiZmZmZmZmqqqqZmZmZmZmIiIiIiIhmZmZ3d3dmZmZmZmZVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3eIiIiIiIiZmZmZmZmqqqq7u7u7u7u7u7u7u7uqqqqqqqqZmZmZmZmZmZmIiIh3d3d3d3d3d3dmZmZmZmZmZmZVVVVVVVVERERVVVVVVVVVVVVERERERERVVVVERERVVVVERERERERERERERERERERVVVVERERVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3eIiIiZmZmZmZmqqqqqqqq7u7vMzMzMzMzMzMy7u7u7u7uqqqqqqqqIiIiIiIiIiIhmZmZmZmZmZmZVVVVERERERERERERERERERERERERERERERERERERERERERERVVVVERERVVVVVVVVmZmZmZmZmZmZmZmZVVVVmZmZVVVVVVVVmZmZmZmZmZmZ3d3eIiIiZmZmqqqqqqqqIiIiIiIhmZmZVVVVVVVVERERERERERERVVVVVVVVmZmZVVVVVVVVmZmZmZmZmZmZ3d3d3d3eIiIiIiIiZmZmZmZmZmZm7u7uqqqrMzMzMzMzMzMzd3d3MzMzMzMzMzMzMzMzMzMy7u7u7u7uZmZl3d3dmZmZVVVVEREREREREREREREQzMzMzMzMzMzNERERERERVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVERERVVVVVVVVVVVVmZmZmZmZ3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3dmZmZmZmZVVVVVVVVVVVVmZmZVVVVmZmZmZmZVVVVmZmZVVVVmZmZmZmZmZmZ3d3dmZmZVVVVEREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREQzMzMzMzMzMzMiIiIREREREREREREiIiIiIiIiIiIREREREREiIiIREREiIiIiIiIiIiIiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIzMzMzMzMiIiIREREREREREREREREiIiIiIiIREREREREiIiIREREREREiIiIREREiIiIREREREREREREiIiIREREiIiIREREREREiIiIREREREREiIiIREREiIiIREREiIiIREREiIiIREREiIiIREREiIiIiIiIREREREREiIiIREREREREiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIREREREREREREiIiIREREiIiIREREREREiIiIiIiIiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIzMzMiIiIiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIREREiIiIiIiIREREREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREiIiIREREREREiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIREREiIiIREREREREiIiIiIiIREREiIiIREREiIiIREREiIiIREREREREREREiIiIREREREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIREREREREiIiIiIiIREREiIiIREREREREiIiIiIiIiIiIREREiIiIiIiIiIiIREREREREiIiIiIiIREREiIiIiIiIREREiIiIREREREREiIiIiIiIzMzMiIiIiIiIiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIzMzMiIiIiIiIzMzMiIiIiIiIiIiIREREREREiIiIREREREREREREiIiIiIiIREREiIiIREREiIiIREREREREiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNERERVVVVVVVVVVVVVVVVmZmZmZmaIiIiIiIiZmZm7u7u7u7vMzMzd3d3u7u7////////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u////////////7u7u////7u7u////////////////7u7u7u7u////7u7u7u7u7u7u3d3d7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d7u7u3d3d3d3d3d3dzMzM3d3d3d3d7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3d7u7u7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3dzMzM3d3dzMzM3d3dzMzMzMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7qqqqqqqqmZmZmZmZqqqqqqqqqqqqqqqqqqqqmZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZqqqqmZmZiIiId3d3iIiId3d3d3d3d3d3ZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3iIiIiIiImZmZmZmZqqqqqqqqu7u7u7u7u7u7qqqqmZmZiIiId3d3d3d3ZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVREREVVVVREREVVVVREREREREREREREREREREREREREREREREVVVVREREVVVVREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmd3d3d3d3d3d3iIiIiIiImZmZmZmZqqqqqqqqqqqqu7u7u7u7zMzMu7u7mZmZiIiIZmZmVVVVVVVVREREREREREREMzMzREREMzMzVVVVREREREREREREREREVVVVVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVZmZmd3d3mZmZqqqqqqqqqqqqmZmZd3d3d3d3ZmZmREREVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3iIiIiIiImZmZqqqqmZmZqqqqqqqqu7u7u7u7zMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7u7u7qqqqmZmZiIiIZmZmVVVVVVVVVVVVREREREREREREMzMzMzMzMzMzREREREREREREVVVVVVVVVVVVREREVVVVVVVVREREREREVVVVREREVVVVZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVREREVVVVZmZmVVVVVVVVVVVVZmZmZmZmmZmZiIiIZmZmZmZmZmZmVVVVREREREREREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiERERIiIiERERIiIiERERIiIiERERIiIiIiIiERERIiIiMzMzIiIiMzMzIiIiIiIiERERIiIiERERERERERERIiIiERERERERIiIiERERERERIiIiERERIiIiERERIiIiERERERERIiIiERERIiIiERERERERIiIiERERERERERERIiIiERERERERERERIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiERERERERERERERERIiIiERERIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERERERIiIiIiIiIiIiIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiERERERERERERIiIiERERIiIiIiIiIiIiIiIiIiIiERERIiIiERERERERIiIiIiIiERERIiIiIiIiMzMzIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERERERIiIiERERIiIiERERERERIiIiERERIiIiIiIiIiIiERERIiIiIiIiERERIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiIiIiIiIiMzMzMzMzIiIiMzMzIiIiIiIiIiIiERERIiIiERERERERIiIiERERIiIiERERERERERERIiIiERERERERERERIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiMzMzMzMzIiIiIiIiERERIiIiIiIiERERERERIiIiERERIiIiIiIiIiIiIiIiERERIiIiIiIiERERERERERERERERIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiERERIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiERERERERIiIiERERERERIiIiIiIiERERIiIiERERIiIiERERIiIiERERIiIiIiIiERERIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREVVVVVVVVVVVVZmZmd3d3d3d3iIiImZmZu7u7zMzM3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7u7u7u7u7u7u7u7u7v///////+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3e7u7t3d3e7u7u7u7t3d3e7u7u7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7t3d3d3d3e7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3e7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3e7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u8zMzMzMzLu7u7u7u7u7u6qqqru7u6qqqqqqqru7u6qqqqqqqpmZmaqqqqqqqru7u6qqqqqqqqqqqpmZmZmZmZmZmZmZmYiIiJmZmZmZmZmZmYiIiHd3d3d3d3d3d2ZmZmZmZnd3d2ZmZnd3d2ZmZlVVVWZmZlVVVWZmZmZmZmZmZlVVVWZmZmZmZlVVVVVVVVVVVWZmZmZmZnd3d3d3d3d3d4iIiJmZmYiIiJmZmZmZmZmZmZmZmZmZmZmZmYiIiHd3d3d3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVURERFVVVURERFVVVURERFVVVURERERERERERERERFVVVVVVVVVVVURERFVVVURERFVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiHd3d4iIiIiIiKqqqru7u6qqqru7u6qqqqqqqoiIiHd3d2ZmZkRERERERERERDMzMzMzM0RERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZlVVVVVVVURERFVVVXd3d4iIiJmZmaqqqpmZmZmZmZmZmXd3d2ZmZmZmZlVVVVVVVVVVVWZmZlVVVWZmZmZmZnd3d3d3d4iIiJmZmaqqqpmZmaqqqqqqqqqqqqqqqszMzLu7u6qqqru7u8zMzMzMzMzMzMzMzMzMzMzMzLu7u6qqqqqqqpmZmXd3d2ZmZmZmZlVVVWZmZlVVVVVVVURERERERERERFVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVURERFVVVVVVVVVVVVVVVURERERERERERERERERERERERFVVVURERERERFVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d1VVVURERERERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIhERESIiIiIiIiIiIiIiIjMzMxERESIiIhERERERERERESIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIhERESIiIhERESIiIhERERERESIiIhERESIiIhERERERESIiIhERERERERERESIiIhERESIiIhERERERESIiIhERERERESIiIhERESIiIhERERERESIiIhERESIiIhERERERESIiIhERERERESIiIhERERERERERERERESIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIhERESIiIhERERERESIiIhERESIiIiIiIjMzMyIiIhERESIiIhERESIiIiIiIiIiIiIiIhERERERERERESIiIhERESIiIhERERERERERESIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIhERERERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIhERESIiIhERESIiIiIiIhERESIiIhERERERESIiIhERERERERERERERERERESIiIjMzMyIiIjMzMzMzMzMzMyIiIiIiIiIiIhERESIiIhERESIiIhERERERERERERERESIiIhERESIiIhERESIiIiIiIiIiIiIiIhERESIiIhERERERERERESIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMyIiIiIiIiIiIhERESIiIhERESIiIhERERERERERESIiIiIiIiIiIhERERERESIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIhERESIiIhERESIiIhERERERESIiIhERERERESIiIhERESIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERFVVVVVVVVVVVWZmZmZmZnd3d4iIiJmZmZmZmaqqqszMzN3d3e7u7u7u7v///////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7////u7u7////u7u7u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7d3d3u7u7d3d3u7u7d3d3u7u7u7u7d3d3u7u7MzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMy7u7vMzMzMzMy7u7u7u7uqqqq7u7u7u7uqqqq7u7u7u7uqqqqqqqqqqqqqqqqqqqq7u7u7u7u7u7vMzMzMzMy7u7u7u7uqqqqqqqqIiIiZmZmZmZmIiIh3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiZmZmIiIiZmZmIiIiIiIiIiIiIiIiIiIhmZmZmZmZVVVVVVVVVVVVVVVVERERERERERERVVVVERERERERERERERERERERERERVVVVERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZ3d3dmZmZmZmaIiIh3d3d3d3eIiIiZmZmZmZmZmZmZmZmIiIiIiIh3d3dVVVVVVVVEREREREQzMzNEREQzMzNEREQzMzNERERERERVVVVERERmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVERERVVVVmZmZ3d3d3d3eIiIiZmZmZmZmZmZmZmZmIiIh3d3dmZmZmZmZmZmZmZmZVVVVmZmZ3d3eIiIiZmZmZmZmZmZmqqqqqqqqZmZmqqqqqqqqqqqqqqqqqqqqZmZmqqqq7u7u7u7vMzMzMzMy7u7u7u7uqqqqqqqqZmZmZmZl3d3dmZmZVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZVVVVmZmZVVVVVVVVVVVVmZmZVVVVVVVVERERERERVVVVVVVVERERVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVEREREREREREQzMzNERERERERVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVEREREREQzMzMzMzMzMzMiIiIzMzMiIiIiIiIzMzMiIiIzMzMzMzMiIiIiIiIiIiIREREiIiIREREREREiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREREREiIiIREREREREiIiIREREiIiIiIiIiIiIREREiIiIiIiIREREiIiIiIiIREREiIiIiIiIREREiIiIREREREREiIiIiIiIiIiIREREREREiIiIREREREREiIiIREREiIiIREREREREREREiIiIREREREREiIiIREREiIiIREREiIiIREREiIiIREREiIiIiIiIREREREREREREiIiIREREiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIiIiIiIiIREREiIiIREREREREiIiIREREREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIREREiIiIiIiIREREREREiIiIREREiIiIREREiIiIiIiIiIiIREREiIiIiIiIREREiIiIiIiIREREiIiIREREiIiIiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIREREiIiIiIiIiIiIREREREREiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIREREREREiIiIREREREREiIiIREREiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIREREiIiIiIiIiIiIREREiIiIiIiIREREREREREREREREiIiIiIiIzMzMzMzMiIiIREREiIiIREREiIiIREREiIiIiIiIzMzMiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMzMzMiIiIiIiIzMzMiIiIzMzMiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIREREiIiIREREREREiIiIREREREREiIiIiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIREREiIiIREREiIiIREREiIiIREREREREREREiIiIiIiIREREzMzMiIiIiIiIREREREREiIiIREREiIiIREREREREiIiIREREREREiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERVVVVVVVVVVVVVVVVVVVV3d3d3d3d3d3d3d3eIiIiIiIiqqqrMzMzMzMzu7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////7u7u////////////////////////////////////////////////////7u7u7u7u7u7u////7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d7u7u7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3dzMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7zMzMu7u7u7u7u7u7u7u7qqqqu7u7qqqqqqqqqqqqqqqqmZmZqqqqu7u7u7u7u7u7u7u7u7u7u7u7zMzMu7u7u7u7mZmZmZmZmZmZmZmZZmZmZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREREREVVVVREREVVVVVVVVVVVVREREVVVVZmZmVVVVVVVVZmZmd3d3ZmZmd3d3d3d3d3d3iIiIiIiImZmZmZmZmZmZmZmZqqqqqqqqmZmZmZmZmZmZd3d3d3d3ZmZmVVVVVVVVREREREREREREREREREREREREREREREREMzMzREREREREREREMzMzREREREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmd3d3iIiIiIiIiIiIiIiIiIiId3d3d3d3VVVVVVVVREREMzMzREREMzMzREREMzMzREREREREREREVVVVVVVVVVVVREREVVVVREREREREVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmiIiImZmZmZmZqqqqmZmZiIiIiIiId3d3ZmZmZmZmZmZmd3d3iIiIiIiImZmZmZmZmZmZmZmZqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqmZmZqqqqu7u7u7u7u7u7u7u7qqqqmZmZmZmZiIiId3d3d3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVZmZmVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVREREREREMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiERERIiIiERERERERIiIiIiIiIiIiIiIiIiIiERERERERIiIiERERIiIiERERERERIiIiERERERERIiIiERERERERIiIiIiIiIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiERERIiIiERERERERIiIiIiIiERERIiIiIiIiIiIiERERIiIiERERIiIiERERERERERERIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiIiIiIiIiERERERERIiIiERERERERIiIiERERIiIiERERIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiERERERERERERIiIiERERERERIiIiERERERERIiIiERERIiIiERERERERIiIiIiIiIiIiIiIiERERIiIiIiIiMzMzIiIiIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERERERERERIiIiIiIiERERERERIiIiIiIiERERIiIiMzMzIiIiERERIiIiERERIiIiERERERERIiIiERERERERIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERERERIiIiERERIiIiERERERERIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiMzMzIiIiIiIiIiIiERERIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERERERERERIiIiIiIiIiIiIiIiERERIiIiERERERERERERIiIiERERERERIiIiERERERERERERIiIiERERIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiMzMzIiIiIiIiMzMzMzMzREREMzMzMzMzMzMzIiIiMzMzREREMzMzREREREREREREREREZmZmVVVVZmZmVVVVVVVVZmZmZmZmVVVVZmZmZmZmiIiIiIiImZmZu7u7zMzMzMzM7u7u////7u7u////////7u7u////////////////7u7u////////////////////////7u7u////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////+7u7t3d3d3d3e7u7u7u7t3d3d3d3d3d3czMzMzMzLu7u7u7u7u7u8zMzMzMzN3d3d3d3d3d3d3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3e7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7v///+7u7u7u7u7u7u7u7t3d3e7u7t3d3e7u7u7u7t3d3e7u7t3d3czMzLu7u6qqqru7u6qqqqqqqqqqqqqqqqqqqqqqqru7u6qqqru7u7u7u6qqqqqqqqqqqqqqqru7u6qqqqqqqqqqqqqqqqqqqqqqqpmZmZmZmZmZmaqqqru7u8zMzLu7u7u7u6qqqpmZmZmZmYiIiGZmZlVVVVVVVVVVVURERERERERERFVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVVVVVURERFVVVURERFVVVVVVVURERFVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d3d3d3d3d5mZmZmZmaqqqqqqqru7u7u7u7u7u7u7u7u7u6qqqpmZmZmZmXd3d3d3d1VVVVVVVURERERERERERERERERERERERERERERERDMzM0RERFVVVURERERERFVVVVVVVURERERERFVVVURERFVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d4iIiIiIiIiIiHd3d2ZmZmZmZlVVVURERERERERERERERERERFVVVVVVVVVVVURERERERERERERERERERERERFVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d3d3d5mZmaqqqqqqqqqqqpmZmZmZmYiIiIiIiIiIiJmZmZmZmZmZmZmZmZmZmaqqqpmZmaqqqqqqqqqqqqqqqqqqqqqqqqqqqpmZmaqqqpmZmaqqqqqqqqqqqqqqqpmZmYiIiHd3d2ZmZnd3d3d3d2ZmZlVVVVVVVURERERERFVVVURERFVVVVVVVURERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZlVVVURERERERFVVVURERFVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVWZmZlVVVURERERERERERERERDMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIiIiIhERESIiIiIiIiIiIiIiIiIiIhERESIiIiIiIhERESIiIhERESIiIiIiIhERESIiIhERERERESIiIiIiIiIiIhERERERESIiIhERESIiIhERESIiIhERERERESIiIhERERERERERESIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIhERERERESIiIhERERERESIiIhERERERESIiIhERERERESIiIhERERERESIiIhERESIiIhERESIiIiIiIiIiIiIiIhERESIiIhERERERESIiIhERESIiIhERERERERERESIiIhERESIiIhERERERESIiIiIiIiIiIhERESIiIhERERERESIiIhERERERESIiIhERESIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIhERESIiIiIiIiIiIhERESIiIhERESIiIhERERERERERERERESIiIiIiIiIiIjMzMyIiIhERESIiIhERESIiIhERERERESIiIiIiIiIiIhERESIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIhERETMzMzMzMyIiIhERERERESIiIhERESIiIhERESIiIiIiIhERESIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIhERERERERERERERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMxERERERESIiIhERESIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIhERESIiIhERESIiIiIiIhERESIiIhERESIiIiIiIiIiIhERESIiIhERESIiIhERESIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM0RERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVXd3d3d3d4iIiKqqqqqqqszMzO7u7u7u7v///////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7////u7u7d3d3d3d3u7u7u7u7d3d3MzMzMzMy7u7uqqqqqqqq7u7u7u7vMzMzMzMzMzMzMzMzd3d3d3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3MzMzd3d3u7u7d3d3u7u7u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7////u7u7////u7u7////////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3u7u7d3d3d3d3MzMzMzMy7u7uqqqqqqqqZmZmqqqqqqqqZmZmqqqqqqqqqqqqqqqqqqqq7u7u7u7uqqqqqqqqZmZmZmZmZmZmqqqqZmZmqqqq7u7uqqqqqqqqqqqqZmZmZmZmZmZmqqqqqqqqqqqq7u7uqqqqqqqqqqqqIiIh3d3dmZmZmZmZVVVVERERERERERERERERERERERERERERERERERERVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVERERVVVVVVVVmZmZmZmZmZmZ3d3eZmZmZmZmqqqqqqqqqqqq7u7uqqqq7u7u7u7uqqqqqqqqqqqqZmZmZmZl3d3dmZmZmZmZmZmZVVVVVVVVERERERERERERERERERERVVVVVVVVERERERERVVVVVVVVERERERERERERERERVVVVERERVVVVERERVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVERERVVVVmZmZ3d3d3d3eIiIiZmZmZmZmIiIiIiIh3d3dmZmZVVVVERERVVVVVVVVERERVVVVVVVVERERVVVVERERERERVVVVERERVVVVERERVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmaIiIiIiIiqqqqqqqq7u7u7u7u7u7uqqqqqqqqZmZmZmZmZmZmZmZmZmZmZmZmZmZmqqqqqqqqqqqqqqqqZmZmqqqqZmZmZmZmZmZmZmZmqqqqZmZmIiIiIiIiIiIhmZmZmZmZmZmZVVVVmZmZ3d3dVVVVERERERERERERERERERERVVVVERERERERERERERERERERERERVVVVERERVVVVVVVVVVVVVVVVmZmZVVVVmZmZ3d3eIiIh3d3dVVVVVVVVmZmZVVVVVVVVVVVVERERVVVVVVVVEREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIiIiIzMzMiIiIzMzMzMzMREREiIiIREREiIiIREREREREREREREREREREREREiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIiIiIiIiIiIiIREREREREiIiIREREREREREREREREiIiIREREREREiIiIREREiIiIREREREREiIiIREREREREiIiIzMzMzMzMiIiIiIiIzMzMiIiIREREiIiIREREREREiIiIREREREREiIiIiIiIiIiIiIiIREREiIiIREREREREiIiIREREiIiIREREREREiIiIREREiIiIiIiIiIiIREREiIiIREREREREiIiIREREREREiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIiIiIiIiIREREiIiIREREiIiIREREiIiIREREREREREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIREREREREiIiIREREiIiIREREREREREREiIiIREREiIiIiIiIiIiIiIiIiIiIREREiIiIREREREREiIiIzMzMiIiIiIiIREREREREiIiIREREiIiIREREiIiIiIiIiIiIREREREREiIiIiIiIREREiIiIiIiIREREiIiIiIiIiIiIzMzMiIiIiIiIREREREREiIiIiIiIREREiIiIREREiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREiIiIiIiIiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIREREiIiIzMzMiIiIiIiIREREREREiIiIREREREREiIiIREREREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREREREREREREREREREiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIREREzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzNERERVVVVVVVVVVVVERERERERERERVVVVmZmZmZmaIiIiIiIiqqqq7u7vMzMzd3d3u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u////7u7u7u7u7u7u7u7u7u7u3d3dzMzMzMzMzMzMzMzMzMzMzMzM3d3d3d3d3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u////7u7u7u7u7u7u7u7u////7u7u////7u7u////7u7u7u7u7u7u7u7u3d3d7u7u3d3d7u7u3d3d7u7u3d3d3d3d3d3d3d3dzMzMu7u7qqqqmZmZmZmZiIiImZmZiIiImZmZmZmZmZmZqqqqqqqqqqqqqqqqqqqqmZmZqqqqiIiIiIiIiIiIiIiImZmZmZmZqqqqqqqqqqqqqqqqqqqqqqqqmZmZqqqqmZmZqqqqqqqqu7u7u7u7u7u7qqqqmZmZmZmZd3d3ZmZmZmZmd3d3ZmZmVVVVREREVVVVVVVVREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVREREVVVVREREVVVVVVVVVVVVZmZmZmZmd3d3d3d3iIiIiIiIiIiIiIiImZmZmZmZqqqqqqqqqqqqqqqqqqqqqqqqmZmZmZmZiIiId3d3d3d3d3d3d3d3ZmZmZmZmVVVVREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVREREVVVVVVVVVVVVREREREREREREVVVVREREVVVVZmZmd3d3iIiImZmZmZmZmZmZiIiIiIiId3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREVVVVREREVVVVVVVVREREVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3qqqqqqqqu7u7zMzMu7u7u7u7mZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZqqqqqqqqmZmZqqqqmZmZmZmZqqqqmZmZmZmZmZmZiIiIiIiId3d3d3d3d3d3VVVVVVVVZmZmZmZmVVVVVVVVREREREREREREMzMzREREMzMzMzMzMzMzMzMzREREMzMzREREREREREREREREREREZmZmZmZmVVVVVVVVZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiERERERERERERIiIiERERIiIiIiIiERERERERIiIiERERIiIiERERERERIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiERERIiIiERERIiIiERERIiIiERERERERIiIiERERERERIiIiERERIiIiMzMzMzMzMzMzIiIiIiIiIiIiERERERERIiIiERERERERIiIiERERIiIiERERERERIiIiIiIiIiIiERERERERERERERERIiIiERERERERIiIiIiIiERERERERERERERERERERIiIiERERERERIiIiERERIiIiERERERERIiIiERERIiIiIiIiERERIiIiIiIiIiIiERERERERIiIiERERERERIiIiERERIiIiERERIiIiIiIiIiIiERERERERIiIiMzMzIiIiIiIiERERIiIiIiIiMzMzMzMzIiIiERERIiIiERERERERERERIiIiERERIiIiIiIiIiIiIiIiERERIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiERERIiIiERERIiIiERERERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiERERIiIiMzMzMzMzIiIiERERERERIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiERERIiIiIiIiIiIiERERIiIiERERIiIiIiIiERERIiIiERERIiIiERERERERIiIiERERIiIiERERMzMzMzMzREREREREIiIiMzMzIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiMzMzIiIiIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiERERIiIiERERERERERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiERERIiIiERERERERIiIiIiIiIiIiERERERERERERIiIiERERERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiERERERERERERIiIiIiIiMzMzIiIiMzMzMzMzIiIiMzMzMzMzREREMzMzIiIiIiIiIiIiMzMzMzMzMzMzREREMzMzREREMzMzREREREREREREREREREREVVVVVVVVREREREREVVVVREREVVVVZmZmZmZmd3d3mZmZmZmZu7u7zMzM3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7t3d3e7u7t3d3d3d3e7u7u7u7u7u7v///+7u7v///////////////////////////////+7u7v///+7u7v///////+7u7v///+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7u7u7t3d3d3d3d3d3d3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7v///+7u7u7u7v///+7u7v///+7u7v///+7u7u7u7u7u7u7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3czMzLu7u6qqqqqqqpmZmYiIiIiIiJmZmZmZmYiIiJmZmZmZmZmZmZmZmZmZmXd3d4iIiIiIiHd3d4iIiIiIiIiIiJmZmaqqqqqqqru7u8zMzLu7u6qqqru7u6qqqqqqqqqqqpmZmZmZmZmZmaqqqqqqqqqqqpmZmZmZmYiIiIiIiIiIiIiIiHd3d3d3d3d3d2ZmZlVVVURERERERERERERERERERERERERERERERERERERERERERERERERERERERERERFVVVWZmZmZmZlVVVWZmZmZmZlVVVVVVVWZmZnd3d4iIiIiIiIiIiIiIiIiIiGZmZnd3d3d3d3d3d4iIiIiIiJmZmZmZmZmZmYiIiHd3d3d3d2ZmZnd3d3d3d4iIiIiIiIiIiHd3d3d3d3d3d1VVVVVVVURERERERERERERERERERDMzMzMzM0RERDMzM0RERDMzM0RERERERERERERERDMzMzMzM0RERDMzM0RERDMzMzMzM0RERFVVVURERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZoiIiIiIiJmZmZmZmaqqqqqqqpmZmZmZmXd3d2ZmZlVVVVVVVVVVVURERERERERERERERERERFVVVURERERERERERERERFVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d4iIiJmZmbu7u7u7u8zMzLu7u7u7u5mZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiHd3d4iIiHd3d3d3d3d3d2ZmZmZmZnd3d2ZmZkRERFVVVVVVVURERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzM0RERFVVVWZmZkRERFVVVWZmZnd3d2ZmZmZmZmZmZmZmZlVVVURERERERERERERERDMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIhERESIiIhERERERERERESIiIhERESIiIhERESIiIhERERERESIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIhERESIiIhERESIiIhERERERESIiIhERESIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERERERESIiIhERESIiIhERERERESIiIhERESIiIhERESIiIhERESIiIhERESIiIhERESIiIhERERERERERESIiIhERESIiIhERESIiIhERESIiIhERESIiIhERESIiIhERESIiIhERERERERERERERESIiIiIiIiIiIiIiIhERERERESIiIhERESIiIhERERERESIiIhERERERESIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIjMzMzMzMxERERERERERERERESIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIhERERERERERERERESIiIiIiIhERESIiIiIiIiIiIiIiIhERESIiIiIiIiIiIkRERDMzMyIiIiIiIiIiIiIiIjMzMyIiIhERERERERERESIiIhERERERERERESIiIhERESIiIiIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIhERESIiIiIiIhERESIiIiIiIiIiIjMzM0RERERERERERCIiIjMzMyIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIhERESIiIiIiIjMzMyIiIhERESIiIhERERERERERESIiIhERERERERERESIiIhERERERERERERERESIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIhERERERERERESIiIhERESIiIhERESIiIhERESIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIhERESIiIhERERERESIiIhERERERESIiIhERERERESIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIhERESIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIjMzM0RERDMzMyIiIiIiIjMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVVVVVURERDMzM0RERERERERERFVVVWZmZlVVVVVVVXd3d3d3d5mZmbu7u8zMzN3d3e7u7u7u7v///////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7u7u7////////////////////////////////u7u7////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3MzMzMzMzMzMzd3d3MzMzd3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7////u7u7////u7u7////////u7u7u7u7////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3MzMzd3d3MzMzMzMzd3d3MzMzMzMzMzMy7u7u7u7u7u7uqqqqZmZmZmZmqqqqqqqqZmZmZmZmIiIiIiIh3d3dmZmZmZmZmZmZmZmZ3d3d3d3eIiIiZmZmqqqq7u7vMzMzMzMzMzMzMzMzMzMzMzMy7u7uqqqqqqqqqqqqZmZmZmZmIiIiZmZmZmZmZmZmqqqqZmZmZmZmZmZmZmZmZmZmZmZmIiIiIiIiIiIh3d3dVVVVVVVVVVVVEREREREQzMzMzMzMzMzNEREQzMzMzMzNERERERERERERERERVVVVVVVVmZmZmZmZmZmZmZmZmZmZ3d3eZmZmqqqqqqqqZmZl3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3eIiIh3d3dmZmZmZmZVVVVVVVVVVVVVVVVmZmZ3d3d3d3d3d3d3d3eIiIh3d3eIiIhmZmZVVVVVVVVVVVVEREREREREREREREREREQzMzMzMzNEREREREQzMzNEREQzMzMzMzNEREQzMzMzMzMzMzNERERERERERERERERERERERERERERVVVVVVVVERERVVVVVVVVmZmZmZmZ3d3d3d3eIiIh3d3eIiIiIiIiqqqqqqqq7u7uqqqqqqqqZmZl3d3dmZmZVVVVEREQzMzMzMzNEREQzMzNEREQzMzNEREQzMzNERERVVVVERERERERVVVVERERVVVVVVVVVVVVmZmZmZmZmZmaIiIh3d3eIiIiqqqq7u7vMzMzMzMy7u7u7u7uZmZmZmZmZmZmIiIiZmZmIiIiZmZmZmZmZmZmIiIiZmZmIiIiIiIiIiIh3d3d3d3d3d3d3d3dmZmZmZmZ3d3eIiIiIiIiIiIhVVVVEREREREREREREREREREREREQzMzNEREREREQzMzNEREREREREREREREREREQzMzNERERVVVVERERERERERERERERERERERERVVVVEREQzMzNEREREREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREREREREREiIiIREREREREREREiIiIREREREREiIiIiIiIREREREREREREREREiIiIREREiIiIREREiIiIREREREREREREREREREREiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREREREREREiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIREREREREREREiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIREREREREREREiIiIiIiIREREiIiIREREREREiIiIREREREREiIiIREREREREREREiIiIiIiIREREREREiIiIREREiIiIiIiIREREiIiIiIiIzMzMiIiIREREiIiIREREiIiIREREiIiIREREREREiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIREREiIiIiIiIREREREREREREiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIREREiIiIiIiIiIiIiIiIREREiIiIREREREREiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIiIiIREREiIiIiIiIREREiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIzMzMzMzMzMzMzMzMiIiIREREiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiJEREQzMzMiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIREREiIiIREREREREREREiIiIiIiIiIiIiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIREREREREiIiIREREiIiIiIiIiIiIiIiIREREiIiIREREiIiIREREREREREREiIiIREREREREREREiIiIiIiIiIiIREREREREiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIREREiIiIREREREREiIiIiIiIzMzMiIiIREREREREiIiIREREiIiIREREiIiIREREiIiIREREzMzMiIiIiIiIREREiIiIiIiIiIiIiIiIREREREREiIiIREREiIiIREREiIiIREREREREiIiIREREREREiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMiIiIzMzMzMzNERERERERVVVVEREREREREREREREREREQzMzNERERERERVVVVVVVVERERVVVVmZmZ3d3eIiIiZmZm7u7vMzMzMzMzd3d3u7u7////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u3d3d3d3d3d3dzMzMu7u7u7u7u7u7zMzM3d3d3d3d3d3d7u7u7u7u7u7u7u7u////7u7u////////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u////7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3dzMzM3d3dzMzMzMzMu7u7zMzM3d3d7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u////7u7u7u7u7u7u////7u7u7u7u////7u7u////7u7u////7u7u////7u7u////7u7u7u7u7u7u7u7u3d3d3d3d3d3dzMzM3d3dzMzM3d3dzMzMzMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7qqqqu7u7qqqqqqqqqqqqmZmZd3d3d3d3ZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiImZmZqqqqqqqqu7u7zMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7u7u7qqqqmZmZiIiIiIiIiIiImZmZmZmZmZmZmZmZqqqqmZmZmZmZmZmZmZmZmZmZmZmZiIiIiIiId3d3ZmZmVVVVVVVVVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVZmZmd3d3iIiImZmZmZmZqqqqiIiIiIiId3d3d3d3d3d3d3d3iIiId3d3iIiImZmZiIiId3d3ZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmVVVVZmZmd3d3d3d3ZmZmZmZmd3d3d3d3d3d3d3d3d3d3ZmZmVVVVVVVVREREREREMzMzREREMzMzREREMzMzREREREREMzMzREREMzMzREREREREREREREREREREREREREREREREREREVVVVZmZmZmZmZmZmiIiIiIiImZmZiIiIiIiIiIiIiIiImZmZiIiImZmZu7u7u7u7u7u7mZmZiIiIZmZmVVVVREREREREMzMzMzMzREREMzMzMzMzMzMzREREREREREREREREVVVVREREREREVVVVVVVVZmZmd3d3d3d3d3d3d3d3d3d3iIiImZmZu7u7u7u7u7u7qqqqmZmZmZmZiIiIiIiIiIiId3d3iIiId3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmd3d3iIiIiIiId3d3ZmZmREREREREZmZmVVVVREREMzMzMzMzREREREREMzMzREREMzMzREREMzMzMzMzMzMzMzMzREREREREMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiMzMzIiIiIiIiERERERERERERERERIiIiERERIiIiERERIiIiIiIiERERERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiIiIiERERERERIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiERERIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiERERERERIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiERERERERERERIiIiIiIiIiIiIiIiERERIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiERERIiIiIiIiIiIiERERIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiMzMzIiIiERERERERERERERERIiIiMzMzIiIiIiIiERERERERIiIiERERERERIiIiIiIiERERERERIiIiIiIiIiIiIiIiERERIiIiMzMzMzMzIiIiERERERERIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiMzMzMzMzMzMzIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiERERIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzIiIiIiIiMzMzMzMzIiIiREREREREMzMzIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiIiIiERERIiIiERERERERIiIiERERIiIiERERERERERERIiIiERERIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiERERERERIiIiERERIiIiERERIiIiIiIiERERIiIiIiIiIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiMzMzIiIiERERERERIiIiERERERERERERIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERERERERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiIiIiMzMzIiIiIiIiMzMzIiIiIiIiIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzREREREREREREMzMzREREVVVVVVVVREREREREREREREREREREVVVVVVVVVVVVZmZmd3d3d3d3d3d3mZmZiIiIqqqq3d3d3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////+7u7u7u7u7u7u7u7szMzMzMzMzMzN3d3czMzN3d3d3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7u7u7u7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3czMzN3d3czMzN3d3e7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7v///+7u7u7u7u7u7v///+7u7v///+7u7v///+7u7v///+7u7v///+7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u7u7u8zMzLu7u7u7u7u7u6qqqqqqqqqqqpmZmaqqqpmZmYiIiGZmZlVVVVVVVVVVVWZmZmZmZnd3d4iIiIiIiIiIiIiIiIiIiKqqqru7u7u7u7u7u8zMzN3d3d3d3czMzN3d3d3d3czMzMzMzMzMzLu7u6qqqpmZmYiIiIiIiIiIiJmZmZmZmaqqqpmZmZmZmaqqqqqqqqqqqpmZmYiIiJmZmYiIiIiIiIiIiHd3d3d3d2ZmZlVVVVVVVURERERERDMzMzMzMzMzM0RERDMzM0RERERERGZmZoiIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiIiIiHd3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiGZmZlVVVVVVVVVVVURERERERERERFVVVURERERERFVVVVVVVVVVVWZmZnd3d3d3d3d3d3d3d5mZmZmZmaqqqpmZmYiIiHd3d2ZmZmZmZlVVVURERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERERERFVVVVVVVWZmZnd3d4iIiJmZmaqqqoiIiIiIiIiIiJmZmYiIiHd3d4iIiIiIiJmZmZmZmaqqqpmZmYiIiHd3d1VVVURERERERERERDMzM0RERDMzMzMzM0RERDMzM0RERERERERERFVVVVVVVVVVVWZmZlVVVXd3d3d3d2ZmZnd3d3d3d3d3d3d3d4iIiIiIiJmZmZmZmZmZmZmZmYiIiHd3d3d3d3d3d2ZmZmZmZnd3d2ZmZnd3d2ZmZnd3d3d3d2ZmZlVVVVVVVVVVVWZmZoiIiJmZmZmZmYiIiHd3d2ZmZmZmZlVVVVVVVURERERERDMzMzMzMzMzMzMzM0RERERERDMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIhERESIiIhERESIiIhERESIiIhERERERERERESIiIiIiIhERESIiIhERESIiIiIiIhERERERESIiIhERERERESIiIhERERERESIiIhERERERESIiIiIiIiIiIhERESIiIhERERERESIiIiIiIhERERERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIhERESIiIiIiIiIiIjMzMzMzMxERESIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERERERERERESIiIhERESIiIiIiIhERERERESIiIhERESIiIhERESIiIhERERERERERESIiIhERESIiIhERESIiIiIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIjMzMzMzMyIiIhERESIiIhERERERERERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIhERERERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIhERERERESIiIhERESIiIhERESIiIiIiIjMzMzMzMyIiIjMzMyIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzM0RERDMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIhERERERESIiIhERESIiIiIiIhERERERESIiIhERERERESIiIhERERERESIiIhERERERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIhERERERESIiIhERERERERERESIiIiIiIhERESIiIhERESIiIhERERERESIiIiIiIiIiIiIiIiIiIhERERERESIiIiIiIiIiIhERESIiIiIiIiIiIhERESIiIhERESIiIhERERERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERERERERERESIiIhERESIiIhERERERESIiIhERESIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERDMzM0RERERERDMzM0RERERERERERERERFVVVWZmZnd3d2ZmZnd3d3d3d3d3d3d3d5mZmaqqqru7u93d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3d3d3MzMzd3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7u7u7u7u7////u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3u7u7d3d3u7u7u7u7////u7u7u7u7u7u7u7u7d3d3u7u7d3d3u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7////u7u7////u7u7////u7u7////u7u7u7u7u7u7d3d3d3d3d3d3d3d3MzMzMzMy7u7u7u7vMzMy7u7u7u7u7u7vMzMy7u7u7u7u7u7uqqqqqqqqqqqqqqqqZmZmZmZmZmZmIiIh3d3eIiIhmZmZmZmZmZmZmZmZVVVV3d3d3d3d3d3eIiIiIiIiIiIiqqqq7u7u7u7vMzMzMzMzMzMzd3d3d3d3d3d3u7u7d3d3d3d3MzMzd3d3MzMy7u7u7u7uqqqqIiIh3d3eIiIiIiIh3d3eIiIiZmZmZmZmqqqqqqqqqqqqZmZmZmZmZmZmIiIiIiIiZmZmZmZmZmZmIiIiIiIhmZmZmZmZVVVVVVVVERERERERERERERERERERVVVV3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3eIiIiIiIh3d3dmZmZERERVVVVERERVVVVERERERERERERERERERERERERERERERERVVVV3d3d3d3d3d3d3d3eIiIiIiIiIiIiZmZmqqqqZmZmqqqqZmZmZmZmIiIhmZmZmZmZEREQzMzNEREQzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNERERERERVVVVmZmZmZmaZmZmZmZmZmZmZmZmIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3eIiIh3d3d3d3eIiIiIiIhmZmZmZmZEREREREREREQzMzMzMzNEREQzMzNERERERERERERERERERERERERERERVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIh3d3dmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVV3d3d3d3eIiIh3d3d3d3dmZmZ3d3eZmZl3d3dEREREREQzMzNEREQzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIzMzMiIiIiIiIREREiIiIiIiIzMzMiIiIREREiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIREREREREiIiIREREiIiIREREiIiIREREiIiIREREzMzMzMzMiIiIREREREREiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIREREiIiIiIiIzMzMiIiIREREiIiIiIiIiIiIiIiIREREiIiIREREiIiIREREREREiIiIiIiIiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIREREiIiIREREiIiIREREiIiIiIiIREREiIiIREREREREiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIREREREREiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREREREiIiIREREiIiIiIiIiIiIzMzMREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIREREiIiIREREiIiIREREiIiIREREREREiIiIiIiIiIiIREREREREiIiIREREREREiIiIREREiIiIiIiIiIiIREREiIiIiIiIiIiIREREREREiIiIREREiIiIREREiIiIREREiIiIREREREREiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREiIiIiIiIiIiIiIiIREREREREiIiIREREiIiIiIiIiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIiIiJEREQzMzNEREQzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIREREiIiIiIiIiIiIiIiIREREiIiIREREiIiIREREREREiIiIREREREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIREREiIiIREREiIiIREREiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIREREiIiIREREiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIREREREREREREREREiIiIiIiIiIiIREREREREiIiIiIiIzMzMiIiIREREREREiIiIiIiIREREiIiIREREiIiIREREREREiIiIREREREREiIiIREREREREiIiIREREiIiIiIiIiIiIzMzMiIiIiIiIiIiIzMzMiIiIzMzMzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzNERERERERERERVVVVmZmZmZmZ3d3eIiIh3d3d3d3eIiIiIiIiIiIiIiIiqqqrMzMzd3d3u7u7////////////////u7u7////////////u7u7////////////////////////////u7u7////////////////////////////////////////////////u7u7////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u3d3dzMzMzMzMzMzMu7u7u7u7zMzM3d3d3d3d7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u7u7u7u7u////7u7u7u7u7u7u3d3d7u7u7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u////7u7u7u7u7u7u7u7uzMzMzMzMzMzMu7u7qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqu7u7qqqqqqqqqqqqu7u7qqqqqqqqqqqqqqqqqqqqqqqqmZmZiIiIiIiIiIiIiIiId3d3d3d3iIiIiIiImZmZiIiImZmZmZmZqqqqu7u7zMzM3d3d3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3du7u7qqqqmZmZiIiId3d3d3d3d3d3ZmZmd3d3d3d3iIiImZmZmZmZiIiImZmZmZmZd3d3iIiIiIiIiIiIiIiIiIiImZmZiIiIiIiIiIiIiIiIZmZmd3d3ZmZmVVVVVVVVVVVVVVVVZmZmiIiId3d3d3d3d3d3d3d3ZmZmd3d3ZmZmZmZmZmZmd3d3ZmZmd3d3d3d3ZmZmREREREREMzMzREREMzMzREREMzMzREREREREREREREREREREVVVVVVVVZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiImZmZmZmZqqqqmZmZmZmZiIiIZmZmZmZmREREREREMzMzREREMzMzREREREREREREREREREREREREVVVVZmZmd3d3mZmZmZmZmZmZiIiImZmZiIiImZmZiIiIiIiIiIiIiIiIiIiId3d3d3d3ZmZmZmZmZmZmZmZmVVVVREREVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3iIiId3d3ZmZmVVVVZmZmVVVVVVVVREREREREREREVVVVREREREREREREREREREREREREREREVVVVREREREREVVVVVVVVd3d3d3d3VVVVREREMzMzMzMzMzMzMzMzMzMzIiIiERERERERIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiMzMzIiIiMzMzIiIiIiIiERERERERERERIiIiIiIiIiIiIiIiERERERERIiIiERERERERIiIiIiIiIiIiIiIiIiIiERERIiIiERERERERERERIiIiERERERERIiIiERERERERIiIiIiIiMzMzIiIiERERERERERERIiIiERERERERIiIiERERIiIiERERERERERERIiIiIiIiIiIiERERERERIiIiIiIiIiIiIiIiERERIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiMzMzMzMzIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERERERIiIiERERIiIiIiIiIiIiERERERERERERERERERERIiIiERERERERIiIiERERIiIiERERERERIiIiIiIiERERIiIiERERIiIiERERERERERERIiIiIiIiIiIiIiIiIiIiIiIiERERERERIiIiERERIiIiERERERERIiIiERERERERIiIiERERIiIiERERIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzMzMzIiIiIiIiERERERERIiIiIiIiERERERERIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiERERERERIiIiERERIiIiIiIiIiIiMzMzIiIiERERERERIiIiERERIiIiERERIiIiERERIiIiIiIiMzMzIiIiIiIiIiIiERERIiIiIiIiIiIiMzMzIiIiIiIiMzMzIiIiIiIiERERERERERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzIiIiERERIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiMzMzIiIiERERERERERERIiIiERERIiIiERERERERIiIiERERIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERERERIiIiERERERERIiIiIiIiERERERERERERIiIiIiIiMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiMzMzIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiERERERERERERERERIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzREREMzMzREREREREREREREREMzMzREREREREVVVVVVVVZmZmd3d3d3d3iIiIiIiIZmZmd3d3iIiImZmZzMzM3d3d7u7u////////////////////////////////////////7u7u////////////////////////////////////////////////////7u7u////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7v///+7u7t3d3d3d3czMzMzMzLu7u8zMzMzMzMzMzN3d3d3d3d3d3e7u7u7u7t3d3e7u7t3d3d3d3d3d3d3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3czMzLu7u6qqqqqqqpmZmYiIiIiIiJmZmYiIiJmZmZmZmZmZmaqqqpmZmZmZmZmZmaqqqpmZmaqqqru7u7u7u6qqqru7u7u7u5mZmaqqqqqqqpmZmZmZmZmZmZmZmaqqqru7u6qqqru7u7u7u7u7u7u7u7u7u8zMzMzMzMzMzN3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3d3d3d3d3czMzLu7u7u7u5mZmYiIiHd3d3d3d3d3d3d3d3d3d2ZmZoiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiJmZmXd3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiHd3d3d3d2ZmZlVVVWZmZlVVVWZmZnd3d2ZmZnd3d2ZmZlVVVURERERERDMzM0RERDMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERGZmZmZmZnd3d4iIiHd3d2ZmZnd3d2ZmZnd3d3d3d2ZmZmZmZlVVVVVVVWZmZnd3d4iIiJmZmZmZmZmZmYiIiHd3d2ZmZmZmZlVVVURERERERERERERERERERFVVVVVVVWZmZmZmZoiIiJmZmZmZmZmZmYiIiJmZmZmZmZmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d2ZmZlVVVURERERERERERERERDMzM0RERDMzMzMzMzMzM0RERDMzM0RERERERDMzM0RERERERERERERERERERFVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d4iIiIiIiHd3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVURERERERERERERERERERERERERERERERDMzMzMzMzMzMyIiIiIiIjMzMyIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIhERERERERERESIiIiIiIhERESIiIhERESIiIiIiIhERESIiIhERESIiIhERERERESIiIhERESIiIhERESIiIiIiIiIiIiIiIhERESIiIhERERERESIiIhERESIiIhERERERESIiIiIiIhERERERESIiIiIiIiIiIhERERERESIiIiIiIiIiIhERESIiIhERESIiIhERESIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIhERESIiIjMzM1VVVURERCIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMyIiIhERESIiIhERESIiIiIiIiIiIjMzMyIiIiIiIhERESIiIhERESIiIhERERERESIiIhERESIiIhERESIiIhERESIiIiIiIhERESIiIhERERERESIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIhERERERESIiIhERESIiIhERESIiIiIiIiIiIjMzMzMzMyIiIiIiIhERESIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIhERESIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIhERERERERERESIiIjMzMyIiIhERERERESIiIhERESIiIhERERERESIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIhERERERERERERERESIiIhERESIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIhERESIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIhERERERESIiIhERETMzMyIiIiIiIhERESIiIhERESIiIhERESIiIhERERERESIiIhERESIiIiIiIhERESIiIiIiIhERESIiIiIiIiIiIhERERERESIiIhERESIiIhERESIiIhERERERESIiIhERESIiIhERESIiIiIiIiIiIhERESIiIiIiIjMzMzMzMyIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIhERESIiIjMzMyIiIhERERERESIiIiIiIhERERERESIiIhERESIiIiIiIiIiIhERESIiIhERESIiIhERESIiIhERERERERERESIiIhERESIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzM0RERERERERERERERERERDMzMzMzM0RERERERFVVVVVVVVVVVWZmZnd3d3d3d3d3d1VVVWZmZnd3d5mZmbu7u93d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////u7u7u7u7u7u7d3d3d3d3MzMzMzMzMzMzMzMzMzMzMzMzd3d3u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7d3d3u7u7u7u7d3d3u7u7d3d3d3d3d3d3MzMy7u7uqqqqZmZmIiIiIiIh3d3eIiIh3d3eIiIiIiIh3d3d3d3eIiIiZmZmIiIiIiIiIiIiZmZmZmZmZmZmZmZmZmZmZmZmZmZmqqqqqqqqqqqqqqqqqqqqZmZmZmZm7u7uqqqq7u7u7u7vMzAD//wAAzN3d3czMzMzMzLu7u6qqqru7u7u7u7u7u8zMzLu7u8zMzMzMzN3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzLu7u5mZmXd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiJmZmZmZmaqqqqqqqqqqqqqqqqqqqpmZmXd3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVURERERERERERDMzM0RERDMzMzMzMzMzMzMzM0RERDMzMzMzM0RERERERGZmZoiIiIiIiJmZmYiIiIiIiIiIiJmZmYiIiHd3d3d3d2ZmZlVVVURERERERERERFVVVVVVVWZmZnd3d4iIiIiIiJmZmYiIiIiIiHd3d3d3d1VVVVVVVURERERERFVVVVVVVWZmZoiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiIiIiHd3d3d3d2ZmZlVVVVVVVTMzMzMzM0RERERERDMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERERERERERERERFVVVVVVVVVVVVVVVURERFVVVVVVVXd3d3d3d5mZmYiIiIiIiHd3d1VVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVURERERERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIhERESIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERERERERERERERESIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERERERERERERERESIiIhERESIiIhERESIiIhERERERESIiIiIiIiIiIiIiIiIiIhERESIiIhERERERESIiIhERESIiIhERERERERERESIiIiIiIhERESIiIiIiIjMzMyIiIhERESIiIhERERERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzM0RERDMzMyIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIhERERERESIiIhERERERESIiIhERESIiIiIiIiIiIhERERERESIiIhERESIiIhERESIiIhERERERESIiIiIiIiIiIiIiIhERERERESIiIhERESIiIhERESIiIiIiIhERESIiIhERESIiIhERERERESIiIhERESIiIhERESIiIhERESIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERERERERERERERESIiIiIiIiIiIiIiIiIiIhERESIiIjMzMyIiIiIiIiIiIhERESIiIiIiIhERESIiIiIiIhERESIiIhERERERESIiIiIiIhERESIiIhERESIiIhERESIiIiIiIjMzMzMzMyIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIhERESIiIhERESIiIhERESIiIiIiIhERESIiIhERESIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERERERERERESIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIiIiIjMzMyIiIhERERERESIiIhERERERESIiIhERESIiIhERERERERERESIiIhERESIiIhERERERESIiIiIiIhERESIiIhERERERERERESIiIhERESIiIhERESIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIjMzMyIiIiIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIhERERERESIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzM0RERERERERERDMzMzMzMyIiIjMzMzMzMzMzM0RERFVVVVVVVVVVVXd3d3d3d1VVVVVVVVVVVWZmZnd3d5mZmbu7u93d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3MzMy7u7vMzMzMzMzMzMzMzMzMzMzd3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7d3d3d3d3d3d27u7uqqqqZmZmIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3eIiIiIiIiIiIh3d3eIiIiIiIiIiIh3d3d3d3d3d3d3d3eIiIiIiIiZmZmqqqqqqqq7u7u7u7u7u7u7u7u7u7u7u7vMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7vMzMzMzMzMzMzd3d3MzMzd3d3d3d3d3d3MzMzMzMyqqqqZmZl3d3eIiIh3d3eIiIiZmZmIiIiZmZmIiIiZmZmZmZmIiIh3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3d3d3d3d3eIiIh3d3eIiIiIiIiIiIiIiIiIiIiZmZmqqqqqqqq7u7u7u7uqqqqqqqqZmZmZmZl3d3d3d3dVVVVVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERVVVWIiIiqqqqqqqqqqqqZmZmZmZmqqqqqqqqZmZmZmZmZmZl3d3dmZmZVVVUzMzNEREQzMzMzMzNERERERERmZmZVVVVmZmZmZmaIiIh3d3eIiIh3d3d3d3d3d3dmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3dmZmZVVVVEREREREQzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzNERERVVVVERERVVVVERERVVVVVVVVmZmZmZmZ3d3eIiIiIiIiZmZmIiIhmZmZVVVVVVVVERERVVVVVVVVVVVVERERERERVVVVEREQzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIREREREREREREiIiIREREREREiIiIiIiIREREiIiIiIiIREREREREiIiIREREiIiIREREREREREREREREREREiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIREREREREiIiIREREiIiIiIiIREREREREiIiIiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIREREREREiIiIREREiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIREREREREiIiIREREREREiIiIiIiIiIiIREREiIiIREREiIiIiIiIREREiIiIiIiIzMzMiIiIzMzMiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIiIiIiIiIiIiIREREiIiIiIiIREREREREiIiIREREiIiIiIiIiIiIREREREREiIiIREREREREiIiIREREREREREREiIiIREREREREiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIREREREREiIiIREREiIiIREREREREiIiIREREiIiIiIiIREREiIiIREREiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIzMzMiIiIREREiIiIiIiIREREiIiIREREiIiIiIiIiIiIREREREREREREiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREREREiIiIREREiIiIREREREREiIiIREREiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIREREiIiIREREiIiIREREiIiIiIiIREREiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMiIiIREREiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREREREiIiIREREREREiIiIiIiIREREREREiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIzMzMiIiIzMzMzMzMiIiIiIiIzMzMzMzMiIiIiIiIzMzMiIiIiIiIREREiIiIiIiIzMzMiIiIREREiIiIiIiIzMzMiIiIREREiIiIREREiIiIREREiIiIREREREREREREiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIzMzMzMzNEREQzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzNERERERERmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmaIiIiqqqrd3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3dzMzMzMzMzMzMu7u7zMzMu7u7zMzMzMzM3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u////7u7u7u7u7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMu7u7qqqqiIiIiIiIiIiId3d3ZmZmd3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3iIiId3d3d3d3iIiIiIiId3d3d3d3ZmZmZmZmd3d3iIiIiIiIiIiImZmZu7u7u7u7u7u7qqqqzMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7zMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM3d3dzMzMu7u7qqqqiIiIiIiId3d3d3d3iIiIiIiImZmZmZmZmZmZmZmZiIiIiIiId3d3d3d3ZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3iIiIiIiImZmZmZmZmZmZmZmZqqqqqqqqmZmZiIiId3d3ZmZmZmZmREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREd3d3iIiImZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZqqqqiIiIZmZmVVVVREREREREREREREREREREREREREREREREREREVVVVVVVVZmZmd3d3iIiIiIiImZmZmZmZmZmZiIiIiIiId3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmd3d3d3d3d3d3ZmZmd3d3VVVVVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREZmZmd3d3d3d3iIiIiIiImZmZmZmZVVVVREREVVVVVVVVREREVVVVREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiERERERERERERIiIiERERIiIiERERIiIiIiIiERERIiIiIiIiERERERERIiIiERERIiIiERERIiIiERERIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiERERIiIiERERERERIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiERERIiIiMzMzMzMzIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiERERERERERERIiIiERERERERIiIiMzMzERERERERERERIiIiIiIiERERIiIiIiIiIiIiERERERERIiIiERERERERIiIiERERERERIiIiIiIiERERERERIiIiERERERERIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiERERIiIiERERERERIiIiERERERERIiIiERERIiIiIiIiERERIiIiERERMzMzMzMzIiIiIiIiMzMzMzMzMzMzIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERERERIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiMzMzMzMzIiIiIiIiMzMzIiIiIiIiERERERERERERIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERERERERERIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiMzMzIiIiIiIiERERIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiERERERERERERIiIiERERIiIiERERIiIiERERERERIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiMzMzIiIiERERIiIiERERERERIiIiERERERERIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzMzMzMzMzMzMzREREREREREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmd3d3qqqqu7u73d3d////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////+7u7u7u7t3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzN3d3d3d3d3d3e7u7u7u7u7u7v///+7u7u7u7v///+7u7v///+7u7v///+7u7u7u7u7u7u7u7u7u7t3d3d3d3czMzMzMzLu7u7u7u6qqqru7u6qqqqqqqoiIiIiIiHd3d3d3d2ZmZmZmZmZmZlVVVXd3d3d3d3d3d3d3d4iIiHd3d4iIiIiIiHd3d3d3d2ZmZnd3d4iIiJmZmZmZmaqqqru7u6qqqpmZmaqqqqqqqru7u7u7u7u7u8zMzMzMzMzMzMzMzLu7u8zMzLu7u7u7u8zMzLu7u7u7u8zMzMzMzMzMzLu7u7u7u8zMzLu7u7u7u7u7u6qqqpmZmYiIiIiIiHd3d3d3d4iIiIiIiIiIiIiIiJmZmYiIiIiIiHd3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVVVVVVVVVWZmZlVVVWZmZmZmZnd3d3d3d2ZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiHd3d4iIiIiIiHd3d2ZmZlVVVVVVVURERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERERERFVVVVVVVWZmZmZmZoiIiIiIiIiIiHd3d3d3d3d3d3d3d4iIiIiIiHd3d2ZmZlVVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERERERFVVVVVVVXd3d4iIiJmZmaqqqpmZmZmZmYiIiHd3d3d3d2ZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZmZmZlVVVURERERERERERERERERERDMzM0RERERERDMzM0RERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVYiIiIiIiHd3d4iIiHd3d1VVVURERFVVVURERERERDMzMzMzMzMzM0RERDMzMzMzMyIiIjMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIhERESIiIiIiIhERESIiIjMzMyIiIiIiIiIiIhERERERESIiIhERESIiIhERESIiIhERESIiIhERESIiIhERERERESIiIhERERERESIiIhERESIiIiIiIiIiIjMzMyIiIiIiIhERESIiIjMzMxERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIhERESIiIhERERERESIiIiIiIhERETMzMzMzMzMzMyIiIhERESIiIhERERERESIiIiIiIiIiIiIiIiIiIjMzMxERESIiIhERESIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIhERESIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIhERESIiIhERERERERERESIiIiIiIiIiIhERERERESIiIhERESIiIhERESIiIhERERERERERESIiIhERESIiIiIiIhERERERESIiIiIiIiIiIiIiIhERERERESIiIiIiIiIiIhERESIiIhERESIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERERERESIiIhERESIiIiIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIhERESIiIhERERERESIiIiIiIiIiIhERERERESIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIhERESIiIiIiIiIiIjMzMzMzMyIiIiIiIhERESIiIhERESIiIhERESIiIhERESIiIiIiIhERESIiIhERESIiIiIiIhERESIiIiIiIhERESIiIhERERERESIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIhERESIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIhERESIiIiIiIhERESIiIiIiIhERESIiIiIiIhERERERESIiIhERESIiIhERESIiIiIiIhERESIiIhERESIiIhERERERERERERERESIiIiIiIiIiIiIiIhERERERESIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIjMzMyIiIhERESIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIjMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzM0RERERERFVVVVVVVVVVVVVVVVVVVURERFVVVXd3d3d3d4iIiKqqqru7u+7u7u7u7v///////////////////////////////////////////////////////////+7u7v///////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////u7u7////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7u7u7u7u7d3d3d3d3d3d3MzMzMzMzMzMzd3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7////u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3MzMzMzMy7u7u7u7u7u7vMzMyqqqqqqqqqqqqqqqqZmZl3d3d3d3dmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3eIiIh3d3d3d3dmZmZmZmZ3d3eIiIiZmZmqqqqqqqqqqqqqqqqqqqqZmZmZmZmZmZmqqqqqqqqqqqqqqqq7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7uqqqq7u7uqqqq7u7uqqqq7u7u7u7uqqqqqqqqZmZmZmZmIiIh3d3d3d3eIiIiIiIiIiIiZmZmIiIiIiIh3d3d3d3dmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZ3d3dmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZVVVVmZmZmZmZVVVVVVVVERERERERERERVVVVVVVVVVVVERERVVVVVVVVmZmZVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVERERERERERERERERVVVVERERERERVVVVERERERERERERERERERERERERERERVVVVmZmZ3d3eIiIiZmZmqqqqqqqqZmZmIiIh3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERERERVVVVVVVVVVVVVVVVEREREREREREREREREREREREQzMzMzMzMzMzNEREQzMzNVVVVVVVVVVVVVVVVVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMiIiIzMzMzMzMiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIREREREREREREiIiIREREiIiIiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIREREiIiIiIiIzMzMzMzMiIiIiIiIiIiIzMzMiIiIREREiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIREREREREiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREREREREREiIiIzMzMiIiIREREiIiIREREREREiIiIREREiIiIzMzMiIiIiIiIzMzMiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzNEREQzMzMzMzMzMzMiIiIREREREREiIiIzMzMzMzMzMzMzMzMREREiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIREREREREREREREREiIiIREREREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIiIiIiIiIzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIREREiIiIREREREREiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIzMzMzMzMREREiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMzMzMREREiIiIREREREREiIiIREREiIiIiIiIREREiIiIREREiIiIiIiIREREiIiIREREiIiIiIiIiIiIREREiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIzMzMREREiIiIiIiIiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMiIiIiIiIREREiIiIiIiIiIiIiIiIREREiIiIREREiIiIzMzMiIiIzMzMiIiIREREREREiIiIREREiIiIREREREREiIiIREREiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIREREiIiIREREiIiIREREREREREREREREiIiIREREiIiIiIiIiIiIzMzMzMzMzMzMzMzNEREQzMzMzMzMiIiIiIiIiIiIiIiIREREiIiIREREREREREREREREiIiIiIiIzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIREREiIiIREREiIiIREREiIiIREREREREiIiIiIiIiIiIREREiIiIiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIREREiIiIiIiIREREREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMzMzNERERERERVVVVVVVVERERERERVVVVVVVV3d3eIiIh3d3eZmZmqqqrd3d3u7u7////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u3d3d3d3d3d3d3d3dzMzM3d3d3d3d7u7u7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3dzMzM3d3du7u7u7u7u7u7zMzMqqqqu7u7qqqqu7u7qqqqqqqqqqqqmZmZiIiIiIiId3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmd3d3iIiImZmZmZmZqqqqqqqqqqqqmZmZmZmZiIiIiIiIiIiIiIiIiIiIiIiImZmZmZmZqqqqmZmZqqqqmZmZmZmZqqqqqqqqqqqqqqqqmZmZmZmZmZmZqqqqqqqqqqqqqqqqu7u7u7u7qqqqmZmZmZmZiIiImZmZmZmZmZmZiIiId3d3d3d3d3d3d3d3ZmZmd3d3ZmZmd3d3ZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmd3d3d3d3VVVVVVVVVVVVREREVVVVREREVVVVVVVVZmZmREREREREREREREREREREMzMzREREREREREREREREREREREREREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVREREVVVVZmZmZmZmd3d3iIiIiIiImZmZmZmZmZmZiIiId3d3ZmZmZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVREREVVVVREREVVVVVVVVREREREREREREREREZmZmd3d3VVVVZmZmd3d3d3d3VVVVREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREMzMzIiIiMzMzIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzREREMzMzIiIiIiIiERERIiIiERERERERERERERERIiIiIiIiERERERERIiIiERERERERIiIiERERERERIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiERERERERIiIiERERIiIiERERERERERERIiIiERERERERIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiERERIiIiIiIiERERIiIiIiIiMzMzIiIiMzMzMzMzMzMzREREMzMzIiIiERERIiIiERERIiIiIiIiMzMzMzMzMzMzMzMzIiIiERERIiIiIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiERERIiIiERERERERIiIiERERERERIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiERERERERERERIiIiERERIiIiERERERERIiIiERERERERIiIiIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiMzMzIiIiERERIiIiMzMzIiIiIiIiIiIiIiIiERERERERIiIiERERIiIiIiIiIiIiERERERERIiIiERERERERIiIiERERERERIiIiIiIiERERIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiIiIiMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiMzMzIiIiERERERERIiIiERERIiIiERERERERIiIiERERIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiERERERERIiIiIiIiIiIiERERERERIiIiIiIiIiIiIiIiIiIiMzMzMzMzREREMzMzMzMzMzMzMzMzIiIiIiIiERERIiIiERERERERERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiERERIiIiERERIiIiERERERERIiIiERERERERERERERERIiIiIiIiIiIiERERIiIiERERERERERERIiIiIiIiERERERERERERIiIiERERIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzREREVVVVVVVVREREVVVVZmZmd3d3d3d3iIiIiIiIiIiIiIiIu7u7zMzM7u7u////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////+7u7v///////////////////////+7u7v///////////////////+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7v///+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7t3d3d3d3d3d3e7u7u7u7u7u7v///+7u7u7u7u7u7t3d3d3d3e7u7t3d3d3d3czMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u6qqqru7u7u7u7u7u7u7u6qqqpmZmZmZmYiIiIiIiHd3d3d3d3d3d2ZmZnd3d2ZmZnd3d3d3d3d3d3d3d5mZmZmZmZmZmYiIiIiIiJmZmYiIiIiIiIiIiJmZmYiIiIiIiJmZmYiIiJmZmYiIiIiIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiJmZmaqqqqqqqru7u7u7u7u7u7u7u6qqqqqqqpmZmYiIiHd3d4iIiIiIiGZmZmZmZnd3d2ZmZmZmZnd3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d4iIiJmZmYiIiJmZmXd3d3d3d1VVVVVVVURERFVVVURERERERERERDMzM0RERDMzM0RERDMzMzMzMzMzMzMzMzMzM0RERDMzM0RERDMzM0RERFVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d3d3d4iIiIiIiIiIiHd3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVURERFVVVURERERERERERERERERERERERERERERERFVVVYiIiIiIiGZmZmZmZpmZmZmZmVVVVVVVVURERERERERERERERDMzM0RERERERERERERERERERDMzMzMzM0RERDMzM0RERDMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIhERESIiIiIiIhERERERESIiIiIiIiIiIhERESIiIiIiIiIiIiIiIhERESIiIiIiIjMzMyIiIiIiIhERERERESIiIhERESIiIhERERERERERESIiIhERERERESIiIhERERERESIiIhERESIiIjMzMyIiIiIiIiIiIhERESIiIiIiIhERESIiIiIiIjMzMzMzMyIiIiIiIhERERERESIiIhERERERESIiIiIiIjMzMzMzMyIiIiIiIhERESIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIhERESIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIhERERERERERESIiIhERERERESIiIhERERERESIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIhERESIiIhERESIiIhERESIiIhERESIiIhERESIiIiIiIhERESIiIhERESIiIhERESIiIhERESIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIhERESIiIiIiIiIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIhERERERERERERERESIiIhERERERESIiIhERESIiIiIiIhERERERESIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMxERESIiIhERESIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIhERESIiIiIiIjMzMyIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIjMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIhERESIiIhERERERESIiIhERERERESIiIiIiIhERESIiIiIiIiIiIiIiIiIiIhERERERESIiIhERESIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIkRERERERDMzMzMzMzMzMyIiIjMzMyIiIhERESIiIiIiIhERERERERERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIiIiIhERESIiIhERESIiIhERESIiIhERESIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIjMzMyIiIjMzMyIiIiIiIjMzMyIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzM0RERERERFVVVVVVVWZmZlVVVWZmZnd3d4iIiHd3d4iIiIiIiKqqqszMzO7u7v///////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3d3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7////u7u7////u7u7////////u7u7////////////////////////////////////////////////////////u7u7u7u7u7u7u7u7u7u7u7u7////u7u7////u7u7u7u7u7u7u7u7d3d3d3d3MzMzMzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7uqqqqqqqq7u7uqqqqqqqqZmZmqqqqZmZmZmZl3d3d3d3dmZmZ3d3d3d3d3d3eIiIiIiIiqqqqqqqqqqqqqqqqZmZmZmZmIiIiIiIiZmZmIiIiIiIiZmZmIiIiIiIiZmZmZmZmIiIiIiIh3d3d3d3dmZmZ3d3dmZmZ3d3d3d3d3d3d3d3eIiIh3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiqqqqqqqqqqqqqqqq7u7uqqqqZmZmZmZmqqqqIiIiIiIh3d3eIiIh3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERERERVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZ3d3eIiIiZmZmqqqqqqqqZmZmIiIiIiIh3d3dmZmZEREREREQzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERERERERERERERERERERERVVVVERERVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVmZmZVVVVVVVVmZmZVVVVVVVVmZmZ3d3dmZmZVVVVVVVVERERVVVVERERVVVVEREREREQzMzNEREQzMzMzMzNERERERERERERERERERERmZmZmZmZmZmZmZmZ3d3d3d3dmZmZEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzMiIiIiIiIiIiIzMzMiIiIzMzMzMzNEREQzMzNEREQzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIREREiIiIREREREREREREiIiIiIiIREREiIiIREREREREiIiIREREREREiIiIREREREREiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIiIiIzMzMiIiIiIiIiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIzMzMzMzMiIiIiIiIREREiIiIREREREREREREREREiIiIiIiIzMzMiIiIREREREREREREiIiIiIiIzMzMiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIzMzMzMzMzMzNEREQzMzMiIiIzMzMzMzMzMzMiIiIREREREREiIiIiIiIiIiIiIiIzMzMzMzMzMzMiIiIiIiIREREREREiIiIiIiIREREiIiIiIiIREREiIiIREREiIiIREREiIiIiIiIzMzMREREREREiIiIzMzMzMzMzMzMREREiIiIREREREREREREiIiIREREiIiIREREREREREREREREiIiIREREREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIREREiIiIREREREREiIiIiIiIREREiIiIREREiIiIREREiIiIREREiIiJEREQzMzMiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIzMzMzMzMzMzNEREREREREREQzMzMzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiJEREQzMzNEREQzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIREREREREiIiIiIiIREREiIiIiIiIREREiIiIiIiIiIiIREREiIiIREREREREREREREREiIiIREREREREREREiIiIREREREREiIiIREREREREiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREREREREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzNERERVVVV3d3dmZmZmZmZ3d3d3d3d3d3eIiIiZmZmqqqrMzMzd3d3u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d7u7u3d3dzMzMzMzMzMzM3d3dzMzMzMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3d3d3d3d3dzMzM3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3dzMzMu7u7zMzMu7u7zMzMzMzMzMzMu7u7zMzMzMzMzMzMu7u7zMzMu7u7qqqqqqqqqqqqqqqqmZmZqqqqqqqqqqqqqqqqmZmZiIiIiIiId3d3iIiImZmZiIiIqqqqqqqqu7u7qqqqqqqqmZmZqqqqmZmZqqqqmZmZmZmZiIiImZmZmZmZmZmZmZmZqqqqiIiIiIiId3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVd3d3d3d3d3d3d3d3iIiIiIiImZmZmZmZmZmZqqqqqqqqqqqqu7u7u7u7qqqqqqqqqqqqqqqqmZmZmZmZd3d3iIiId3d3d3d3ZmZmZmZmZmZmZmZmVVVVVVVVREREVVVVREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmd3d3iIiImZmZmZmZmZmZmZmZiIiId3d3VVVVREREREREREREREREMzMzREREMzMzREREREREREREMzMzREREREREREREMzMzREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREVVVVVVVVVVVVVVVVVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiMzMzMzMzMzMzMzMzERERIiIiIiIiIiIiIiIiERERERERIiIiERERERERIiIiERERIiIiERERERERIiIiERERIiIiIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiERERIiIiERERERERIiIiERERERERERERERERIiIiMzMzIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiMzMzIiIiIiIiERERIiIiERERERERERERIiIiIiIiMzMzMzMzMzMzIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiERERIiIiIiIiMzMzIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiMzMzMzMzIiIiIiIiIiIiERERIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiMzMzIiIiIiIiERERIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiERERIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiERERERERIiIiERERIiIiERERIiIiERERIiIiIiIiERERERERIiIiERERIiIiIiIiERERIiIiREREMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiERERERERIiIiERERERERIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzREREMzMzREREMzMzMzMzIiIiERERERERERERIiIiERERIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERERERIiIiERERERERIiIiIiIiIiIiMzMzMzMzMzMzIiIiERERIiIiIiIiMzMzIiIiIiIiERERIiIiIiIiIiIiMzMzIiIiMzMzIiIiREREREREVVVVMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiERERERERIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiERERIiIiMzMzIiIiIiIiIiIiIiIiERERIiIiIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERERERIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiREREVVVVd3d3ZmZmVVVVZmZmd3d3iIiIiIiImZmZqqqqu7u73d3d7u7u7u7u////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7u7u7t3d3e7u7t3d3d3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3czMzMzMzN3d3czMzMzMzN3d3czMzN3d3d3d3e7u7t3d3e7u7u7u7t3d3d3d3d3d3e7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3czMzMzMzLu7u7u7u7u7u7u7u8zMzMzMzMzMzMzMzMzMzN3d3d3d3e7u7u7u7u7u7t3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzLu7u7u7u5mZmaqqqqqqqqqqqqqqqru7u7u7u7u7u7u7u7u7u7u7u8zMzLu7u7u7u6qqqqqqqqqqqpmZmaqqqqqqqqqqqpmZmaqqqpmZmZmZmZmZmZmZmZmZmaqqqru7u7u7u6qqqqqqqqqqqqqqqpmZmYiIiJmZmZmZmZmZmZmZmZmZmYiIiJmZmZmZmZmZmYiIiHd3d2ZmZmZmZlVVVVVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d2ZmZmZmZnd3d3d3d4iIiIiIiKqqqqqqqqqqqqqqqru7u7u7u7u7u7u7u8zMzLu7u7u7u7u7u6qqqpmZmZmZmYiIiIiIiIiIiHd3d2ZmZmZmZlVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERERERERERFVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVURERFVVVVVVVWZmZnd3d5mZmZmZmYiIiHd3d4iIiIiIiGZmZmZmZlVVVURERDMzM0RERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERERERERERGZmZlVVVURERERERDMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERERERFVVVURERFVVVVVVVVVVVVVVVWZmZkRERERERDMzMzMzMyIiIiIiIjMzMzMzMzMzMyIiIiIiIjMzMzMzM0RERDMzMzMzMyIiIjMzMyIiIjMzMyIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzMyIiIiIiIhERERERESIiIiIiIiIiIiIiIhERERERESIiIhERERERESIiIiIiIhERESIiIhERESIiIiIiIiIiIhERESIiIhERESIiIhERERERESIiIhERESIiIhERESIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIhERESIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERERERERERERERERERESIiIjMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIhERERERERERESIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMyIiIjMzMzMzMzMzMyIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIhERESIiIhERESIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIhERESIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIjMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIhERESIiIiIiIiIiIhERESIiIiIiIhERERERESIiIhERESIiIhERERERESIiIiIiIhERESIiIiIiIiIiIiIiIiIiIjMzMzMzM0RERERERDMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzM0RERDMzMzMzMyIiIiIiIhERESIiIhERESIiIhERESIiIhERESIiIhERESIiIiIiIhERERERERERERERESIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzM1VVVURERERERDMzMzMzMzMzMyIiIiIiIiIiIiIiIhERESIiIiIiIhERERERESIiIhERESIiIhERESIiIhERERERESIiIiIiIhERESIiIhERERERERERESIiIhERESIiIhERERERESIiIhERESIiIhERESIiIhERESIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIhERERERESIiIhERESIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIiIiIhERESIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMyIiIjMzM1VVVVVVVURERERERFVVVWZmZnd3d4iIiIiIiJmZmZmZmbu7u93d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7////u7u7u7u7u7u7d3d3d3d3d3d3d3d3MzMzMzMzMzMzd3d3d3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMzMzMyqqqqqqqqZmZmZmZmZmZmqqqqqqqqqqqq7u7uqqqq7u7uqqqq7u7uqqqqqqqqqqqqZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmqqqqZmZmZmZmqqqqqqqqqqqq7u7u7u7u7u7u7u7u7u7uqqqqqqqqZmZmZmZmqqqqZmZmZmZmIiIiZmZmZmZmZmZmIiIiIiIh3d3dmZmZVVVVVVVVVVVVERERERERERERERERVVVVERERVVVVERERERERVVVVVVVVmZmZ3d3dmZmZmZmZ3d3eIiIiZmZmqqqqqqqq7u7vMzMzMzMzd3d3MzMzd3d3MzMzMzMzMzMzMzMy7u7u7u7uqqqqqqqqqqqqZmZmIiIh3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERERERERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVmZmZVVVVVVVVVVVVVVVVERERERERVVVVERERERERERERERERERERVVVVmZmZVVVVmZmZmZmZ3d3d3d3eIiIiIiIh3d3dmZmZmZmZmZmZVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERVVVVERERVVVVVVVVmZmZVVVVmZmZVVVVVVVVVVVVVVVVERERERERVVVVmZmZ3d3dmZmZVVVVEREQzMzMzMzMzMzMzMzMzMzNERERERERERERERERERERERERVVVVVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMiIiIzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMiIiIiIiIzMzMzMzMiIiIiIiIzMzMiIiIiIiIREREREREiIiIiIiIREREREREREREiIiIREREREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREREREREREiIiIREREiIiIREREiIiIREREREREiIiIREREREREREREiIiIREREREREREREiIiIiIiIzMzMREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIREREiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIREREREREiIiIiIiIREREiIiIREREzMzMiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIREREREREiIiIREREiIiIiIiIREREiIiIiIiIzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMiIiIzMzMiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREREREiIiIiIiIREREREREiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzMiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMREREREREiIiIiIiIiIiIiIiIREREREREiIiIREREiIiIREREiIiIiIiIREREiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIREREiIiIREREiIiIREREREREREREREREiIiIREREREREiIiIREREiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiJEREREREREREQzMzMzMzMiIiIiIiIiIiIzMzMiIiIiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIREREREREiIiIREREiIiIiIiIREREiIiIREREiIiIREREREREREREiIiIREREiIiIREREREREREREiIiIREREREREiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREREREiIiIREREiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIREREiIiIREREiIiIiIiIiIiIzMzMiIiIzMzMzMzMiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERVVVVmZmZmZmZ3d3eIiIiIiIiIiIi7u7vMzMzu7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3d3d3d7u7u3d3d3d3d3d3d7u7u7u7u7u7u3d3d7u7u3d3d3d3d7u7u3d3d3d3d7u7u7u7u7u7u7u7u////////////////////7u7u7u7u////////7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d7u7u7u7u7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3dzMzMu7u7qqqqqqqqqqqqqqqqqqqqmZmZqqqqqqqqqqqqqqqqmZmZmZmZqqqqmZmZmZmZmZmZiIiId3d3d3d3iIiImZmZmZmZqqqqmZmZmZmZmZmZqqqqmZmZqqqqqqqqu7u7u7u7u7u7u7u7zMzMzMzMu7u7u7u7u7u7qqqqqqqqmZmZmZmZmZmZiIiId3d3ZmZmVVVVVVVVVVVVREREREREREREREREMzMzREREREREREREREREREREVVVVVVVVZmZmZmZmd3d3d3d3d3d3iIiIiIiImZmZqqqqu7u7u7u7zMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMu7u7u7u7qqqqqqqqiIiIiIiIiIiId3d3d3d3ZmZmZmZmZmZmVVVVVVVVREREVVVVREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREVVVVVVVVREREREREVVVVREREREREREREREREREREVVVVREREVVVVVVVVVVVVZmZmd3d3ZmZmZmZmZmZmd3d3iIiIZmZmVVVVREREREREREREMzMzMzMzREREREREMzMzREREREREREREREREREREREREREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVZmZmVVVVZmZmiIiImZmZVVVVREREREREMzMzREREREREMzMzMzMzMzMzREREREREREREREREREREREREMzMzMzMzMzMzMzMzIiIiIiIiMzMzMzMzMzMzREREMzMzMzMzREREMzMzMzMzIiIiIiIiIiIiIiIiMzMzMzMzREREREREREREMzMzMzMzIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiERERIiIiIiIiIiIiERERIiIiERERERERIiIiERERERERIiIiERERERERIiIiERERIiIiERERERERIiIiERERIiIiMzMzIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERERERERERERERIiIiMzMzIiIiERERERERERERERERIiIiIiIiERERERERIiIiIiIiIiIiIiIiERERIiIiERERERERERERIiIiIiIiIiIiMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzIiIiMzMzIiIiMzMzIiIiIiIiMzMzIiIiMzMzMzMzIiIiMzMzIiIiIiIiERERIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERERERERERIiIiERERERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiMzMzIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzMzMzREREMzMzMzMzMzMzMzMzIiIiERERERERIiIiIiIiIiIiIiIiERERIiIiERERERERERERIiIiIiIiIiIiERERIiIiIiIiMzMzMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzIiIiMzMzIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiERERERERIiIiERERERERERERIiIiIiIiERERIiIiERERIiIiERERIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERERERIiIiIiIiMzMzIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiMzMzERERIiIiIiIiMzMzIiIiIiIiREREMzMzMzMzMzMzMzMzIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERERERERERERERIiIiERERIiIiERERERERERERIiIiERERIiIiERERERERIiIiERERIiIiIiIiIiIiIiIiIiIiERERERERIiIiERERIiIiERERERERIiIiERERERERERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREZmZmZmZmd3d3d3d3ZmZmiIiImZmZqqqqzMzM3d3d7u7u////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7t3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzN3d3czMzMzMzMzMzMzMzN3d3d3d3d3d3d3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7u7u7u7u7t3d3e7u7t3d3e7u7t3d3e7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7v///+7u7u7u7u7u7u7u7u7u7v///+7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3czMzLu7u6qqqqqqqqqqqqqqqpmZmZmZmZmZmZmZmZmZmZmZmaqqqoiIiJmZmYiIiIiIiHd3d2ZmZnd3d3d3d4iIiKqqqoiIiIiIiHd3d4iIiIiIiIiIiJmZmZmZmZmZmZmZmaqqqqqqqru7u7u7u7u7u7u7u7u7u8zMzKqqqqqqqqqqqpmZmYiIiIiIiHd3d1VVVVVVVVVVVURERFVVVURERDMzMzMzM0RERDMzM0RERERERERERFVVVVVVVVVVVWZmZmZmZnd3d4iIiHd3d4iIiJmZmaqqqru7u7u7u7u7u8zMzMzMzMzMzMzMzMzMzMzMzMzMzN3d3d3d3czMzMzMzLu7u7u7u5mZmZmZmZmZmYiIiIiIiIiIiIiIiHd3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERFVVVURERFVVVURERERERERERFVVVURERERERERERERERFVVVVVVVWZmZlVVVVVVVWZmZmZmZlVVVVVVVXd3d3d3d3d3d1VVVVVVVURERFVVVVVVVURERERERERERDMzMzMzMzMzMzMzM0RERERERERERERERERERERERERERFVVVURERFVVVVVVVVVVVWZmZoiIiHd3d1VVVXd3d5mZmXd3d1VVVURERDMzM0RERERERERERDMzMzMzMzMzM0RERERERDMzM0RERDMzMzMzMyIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzM0RERERERERERERERDMzMyIiIjMzMyIiIjMzMzMzMzMzM0RERDMzM0RERERERDMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIhERESIiIiIiIiIiIhERERERESIiIhERERERESIiIhERESIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIhERESIiIhERESIiIiIiIhERESIiIhERESIiIiIiIjMzMyIiIhERESIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIjMzM0RERERERFVVVTMzMzMzM0RERDMzMzMzMyIiIjMzMyIiIiIiIjMzMyIiIjMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIhERERERESIiIhERESIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIhERESIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIiIiIjMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMyIiIjMzMyIiIhERESIiIiIiIiIiIiIiIhERESIiIhERESIiIhERESIiIhERESIiIiIiIjMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMyIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzM0RERDMzM0RERDMzMyIiIjMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzMyIiIjMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzMzMzMyIiIiIiIhERESIiIhERERERESIiIhERERERESIiIhERERERESIiIiIiIhERESIiIiIiIkRERDMzMyIiIiIiIiIiIhERESIiIhERESIiIhERESIiIiIiIiIiIjMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIjMzMyIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIhERESIiIhERESIiIhERESIiIhERERERESIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIhERESIiIjMzMyIiIiIiIiIiIhERERERESIiIhERESIiIhERERERESIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIhERESIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERERERERERFVVVVVVVWZmZnd3d2ZmZnd3d5mZmaqqqru7u8zMzO7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3MzMzd3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7////u7u7////u7u7////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d27u7uqqqqqqqqqqqqZmZmZmZmZmZmZmZmZmZmZmZmqqqqqqqqZmZmIiIiIiIh3d3d3d3dmZmZmZmZmZmZ3d3eIiIiIiIh3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiZmZmZmZmZmZmZmZmqqqq7u7uqqqqqqqq7u7u7u7u7u7uqqqqqqqqIiIiIiIh3d3dmZmZVVVVVVVVVVVVEREREREREREREREQzMzNERERERERERERERERERERERERVVVVVVVVmZmZmZmZmZmZmZmZ3d3eIiIiqqqq7u7vMzMzMzMzMzMzMzMy7u7u7u7u7u7vMzMzMzMzMzMzMzMzMzMzMzMy7u7u7u7uqqqqZmZmIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3dmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVERERERERVVVVERERERERVVVVEREREREQzMzNEREREREREREREREQzMzNERERERERERERVVVVVVVVmZmZVVVVmZmZmZmZVVVVVVVVVVVVmZmZmZmZVVVVVVVVERERERERERERVVVVEREREREQzMzMiIiIzMzMzMzNEREREREREREREREQzMzNERERERERERERERERERERVVVVVVVVERERmZmZ3d3dmZmZmZmaZmZl3d3dVVVVEREQzMzMzMzNEREREREQzMzMzMzNEREQzMzNEREQzMzMiIiIzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIzMzMzMzNEREREREREREQzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMiIiIiIiIiIiIiIiIzMzMzMzMREREREREREREiIiIiIiIREREREREiIiIiIiIzMzMiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIREREiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIiIiIiIiIREREREREREREiIiIREREiIiIiIiIREREREREiIiIzMzMiIiIiIiIiIiIiIiIREREREREiIiIiIiIREREiIiIiIiIiIiIiIiIzMzMzMzMzMzNEREQzMzMzMzNEREREREQzMzMzMzMiIiIzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzMiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIREREiIiIREREiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIREREREREiIiIREREREREiIiIREREREREiIiIiIiIzMzMiIiIiIiIiIiIREREREREREREiIiIiIiIiIiIzMzMREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIREREREREiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzMzMzMzMzMiIiIzMzMzMzNEREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzMiIiIzMzMzMzMiIiIiIiIiIiIzMzMiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMiIiIzMzMzMzNEREQzMzMzMzMiIiIiIiIREREiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIREREREREiIiIzMzMzMzMiIiIiIiIiIiIREREREREiIiIREREREREiIiIiIiIzMzMiIiIzMzMzMzMiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiJEREQzMzMzMzMiIiIiIiIzMzMiIiIREREREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREREREiIiIREREREREiIiIREREREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIREREiIiIiIiIREREiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERVVVVVVVVmZmZ3d3d3d3eIiIiqqqqqqqq7u7vu7u7u7u7////////u7u7////////////////u7u7////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u3d3dzMzMzMzMzMzMzMzM3d3dzMzMzMzMzMzMzMzM3d3dzMzM3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u3d3d7u7u3d3d3d3d7u7u3d3d7u7u3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u////7u7u7u7u7u7u////7u7u7u7u////7u7u////7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMu7u7qqqqqqqqqqqqmZmZmZmZmZmZqqqqqqqqmZmZiIiImZmZiIiId3d3d3d3ZmZmd3d3d3d3VVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3iIiId3d3d3d3d3d3iIiId3d3iIiImZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZiIiImZmZiIiId3d3ZmZmZmZmZmZmZmZmZmZmVVVVREREREREVVVVREREREREREREVVVVREREVVVVREREVVVVVVVVZmZmZmZmd3d3iIiIqqqqu7u7zMzMzMzMu7u7u7u7zMzMu7u7u7u7u7u7u7u7zMzMzMzMzMzMzMzMu7u7u7u7mZmZmZmZiIiId3d3ZmZmd3d3ZmZmd3d3iIiId3d3iIiIiIiIiIiIiIiIiIiIiIiId3d3iIiIiIiIiIiId3d3d3d3ZmZmd3d3VVVVVVVVVVVVREREVVVVVVVVREREVVVVVVVVREREREREREREMzMzREREMzMzREREREREREREREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVZmZmZmZmVVVVVVVVREREVVVVVVVVREREREREREREMzMzIiIiIiIiMzMzMzMzMzMzREREREREREREMzMzMzMzMzMzREREREREREREREREVVVVREREREREVVVVZmZmVVVVd3d3VVVVREREMzMzMzMzMzMzREREREREREREMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiMzMzIiIiIiIiIiIiMzMzMzMzREREMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzREREMzMzMzMzMzMzIiIiERERERERERERIiIiIiIiIiIiIiIiERERIiIiERERERERERERIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzIiIiERERIiIiERERIiIiIiIiIiIiIiIiERERERERIiIiERERIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiMzMzMzMzIiIiMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzIiIiIiIiERERERERIiIiERERIiIiERERERERIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzREREMzMzMzMzMzMzMzMzREREMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiMzMzMzMzIiIiIiIiMzMzMzMzIiIiMzMzREREREREIiIiIiIiIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzIiIiERERIiIiIiIiIiIiMzMzMzMzIiIiIiIiERERIiIiERERIiIiERERIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREREREREREREREMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzREREREREMzMzIiIiIiIiIiIiERERERERIiIiERERERERIiIiERERERERERERERERIiIiERERIiIiIiIiMzMzIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzREREREREMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiMzMzMzMzIiIiIiIiERERERERIiIiIiIiIiIiERERIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzIiIiERERERERERERIiIiIiIiERERIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiMzMzIiIiERERIiIiIiIiIiIiERERERERIiIiERERIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzREREMzMzIiIiMzMzMzMzMzMzREREREREREREVVVVZmZmZmZmZmZmd3d3mZmZmZmZmZmZzMzM7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///93d3czMzMzMzMzMzLu7u8zMzN3d3czMzN3d3czMzMzMzN3d3d3d3e7u7t3d3e7u7t3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7u7u7u7u7u7u7u7u7v///+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7v///+7u7u7u7u7u7u7u7t3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzLu7u6qqqqqqqqqqqqqqqqqqqru7u6qqqoiIiIiIiIiIiGZmZmZmZlVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiIiIiJmZmZmZmZmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d2ZmZlVVVWZmZlVVVVVVVURERFVVVURERFVVVVVVVVVVVWZmZnd3d3d3d4iIiJmZmaqqqqqqqru7u6qqqru7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqoiIiIiIiHd3d3d3d3d3d2ZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiJmZmZmZmaqqqqqqqqqqqpmZmZmZmYiIiHd3d2ZmZmZmZlVVVVVVVVVVVURERERERERERERERERERERERERERERERERERERERERERFVVVURERFVVVVVVVWZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVVVVVVVVVVVVVTMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzM0RERERERDMzMzMzMzMzM0RERERERERERERERFVVVVVVVURERERERFVVVVVVVVVVVURERDMzMzMzMyIiIjMzMzMzMzMzM0RERDMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIjMzMzMzMzMzMyIiIjMzMzMzMyIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMyIiIiIiIiIiIhERESIiIjMzMyIiIhERESIiIhERESIiIhERESIiIiIiIjMzMyIiIiIiIhERERERESIiIhERERERESIiIhERESIiIiIiIiIiIiIiIhERESIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIhERESIiIiIiIjMzMyIiIiIiIjMzMzMzMzMzM0RERDMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMyIiIhERERERESIiIhERERERERERERERESIiIhERERERESIiIhERESIiIiIiIjMzMzMzMyIiIjMzMyIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIjMzMyIiIjMzM0RERDMzMyIiIjMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMyIiIiIiIhERERERESIiIiIiIjMzMyIiIiIiIhERESIiIiIiIiIiIiIiIhERERERESIiIhERESIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMyIiIjMzMyIiIjMzM1VVVURERCIiIiIiIiIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMyIiIiIiIjMzMyIiIiIiIhERESIiIjMzMyIiIjMzMzMzMyIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzM0RERDMzM0RERERERDMzM0RERFVVVVVVVURERERERERERDMzMzMzMyIiIjMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzMyIiIiIiIhERERERESIiIhERERERESIiIhERERERESIiIiIiIhERERERESIiIhERERERESIiIjMzMyIiIhERESIiIhERESIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIjMzMyIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzM1VVVURERDMzMyIiIiIiIiIiIiIiIhERERERESIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERERERESIiIhERESIiIhERERERESIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIhERESIiIhERESIiIhERESIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIjMzMyIiIiIiIjMzMyIiIiIiIhERESIiIhERERERESIiIhERESIiIjMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzM0RERERERFVVVURERFVVVWZmZmZmZoiIiIiIiKqqqszMzN3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////u7u7u7u7MzMzMzMzMzMzMzMzd3d3MzMzd3d3d3d3d3d3d3d3d3d3u7u7d3d3d3d3u7u7d3d3d3d3MzMzMzMzMzMzd3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7u7u7d3d3u7u7u7u7u7u7u7u7////////u7u7////////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3MzMzd3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3MzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7uZmZmZmZmIiIh3d3dVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3eIiIh3d3d3d3eIiIiIiIh3d3eIiIh3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIiZmZmIiIiIiIh3d3eIiIh3d3d3d3eIiIiIiIh3d3dmZmZmZmZmZmZmZmZVVVVmZmZVVVVmZmZ3d3eIiIiZmZmqqqqZmZmZmZmZmZmZmZmqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqq7u7uqqqqZmZmIiIiIiIh3d3d3d3d3d3dmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZ3d3eIiIiIiIiIiIiZmZmZmZmZmZmqqqqqqqqqqqqqqqq7u7uqqqqqqqqZmZmIiIiIiIhmZmZmZmZVVVVVVVVERERERERERERERERERERERERERERERERVVVVERERERERVVVVVVVVmZmZmZmZ3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZERERERERERERERERERERVVVVEREQzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzNERERERERERERVVVVEREREREREREREREREREQzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIREREiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREREREREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIREREiIiIiIiIiIiIREREiIiIiIiIiIiIREREiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMiIiIiIiIREREiIiIREREiIiIiIiIiIiIREREREREiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIzMzMiIiIzMzMiIiIzMzMzMzMiIiIiIiIzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIzMzMzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIREREREREiIiIiIiIzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIREREiIiIzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIiIiIREREiIiIiIiIiIiIzMzMzMzMiIiIiIiIREREiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIREREiIiIzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzNEREQzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMiIiIzMzMzMzMREREiIiIiIiIiIiIzMzMzMzMzMzMzMzMiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzNEREQzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREREREQzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMiIiIzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREREREQiIiIREREREREiIiIREREiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIzMzMiIiIiIiIiIiIiIiJERERVVVUzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIzMzMiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIREREiIiIREREREREiIiIREREREREiIiIREREiIiIiIiIiIiIiIiIzMzMiIiIiIiIzMzMiIiIzMzMzMzMiIiIREREREREiIiIiIiIREREiIiIiIiIzMzMiIiIiIiIzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIREREREREiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIzMzNEREQzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzNERERERERVVVVVVVVmZmZ3d3eIiIiZmZmqqqq7u7vMzMzu7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u3d3d7u7u7u7u7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzM3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u////7u7u7u7u7u7u////7u7u////7u7u////7u7u////7u7u7u7u7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzMzMzMzMzMzMzMu7u7u7u7zMzMzMzMzMzMzMzMzMzM3d3dzMzMzMzMzMzMzMzMu7u7qqqqqqqqmZmZd3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZiIiIiIiIiIiIiIiId3d3d3d3d3d3iIiImZmZmZmZmZmZmZmZiIiImZmZmZmZiIiImZmZiIiImZmZmZmZmZmZmZmZmZmZmZmZmZmZiIiIiIiIZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3iIiImZmZqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqmZmZmZmZiIiIiIiId3d3ZmZmVVVVREREREREREREMzMzMzMzREREREREREREREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmVVVVREREREREREREVVVVZmZmZmZmd3d3VVVVREREMzMzMzMzMzMzMzMzREREMzMzREREREREREREMzMzREREREREREREMzMzREREMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzIiIiERERERERIiIiMzMzIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiERERIiIiIiIiMzMzIiIiIiIiERERIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiERERIiIiERERERERERERIiIiIiIiERERIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREREREMzMzIiIiIiIiIiIiERERERERIiIiIiIiIiIiERERERERIiIiERERERERIiIiIiIiIiIiIiIiERERIiIiMzMzIiIiERERIiIiERERIiIiIiIiIiIiIiIiMzMzIiIiIiIiMzMzMzMzMzMzIiIiMzMzMzMzREREMzMzIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiERERIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiMzMzIiIiIiIiERERIiIiMzMzIiIiMzMzIiIiIiIiERERERERERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzIiIiIiIiMzMzMzMzIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzIiIiERERIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzREREREREREREMzMzREREMzMzREREMzMzMzMzMzMzREREVVVVREREREREREREMzMzREREMzMzMzMzMzMzREREREREMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREMzMzIiIiIiIiERERIiIiERERERERIiIiERERERERERERIiIiERERERERIiIiIiIiERERERERIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiREREREREMzMzIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiERERIiIiERERIiIiERERERERIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiERERERERIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiREREMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREREREVVVVVVVVZmZmd3d3iIiIiIiIiIiIqqqqzMzM3d3d7u7u7u7u////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7u7u7u7u7u7u7v///+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7u7u7u7u7t3d3e7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7v///+7u7v///+7u7v///+7u7v///+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3czMzMzMzLu7u8zMzMzMzMzMzMzMzMzMzLu7u6qqqqqqqru7u6qqqru7u8zMzMzMzLu7u8zMzMzMzMzMzN3d3czMzLu7u6qqqpmZmYiIiIiIiHd3d2ZmZmZmZnd3d2ZmZmZmZlVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVWZmZmZmZlVVVWZmZmZmZmZmZnd3d3d3d3d3d4iIiIiIiIiIiHd3d4iIiIiIiIiIiIiIiIiIiJmZmYiIiIiIiJmZmZmZmYiIiJmZmZmZmZmZmaqqqpmZmZmZmZmZmZmZmZmZmZmZmYiIiJmZmYiIiJmZmZmZmYiIiJmZmZmZmZmZmYiIiGZmZmZmZlVVVWZmZlVVVWZmZlVVVVVVVWZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiIiIiIiIiJmZmaqqqpmZmZmZmaqqqpmZmaqqqqqqqpmZmZmZmZmZmZmZmZmZmYiIiJmZmYiIiHd3d2ZmZmZmZlVVVURERERERERERERERERERFVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVWZmZmZmZlVVVVVVVVVVVWZmZmZmZlVVVWZmZoiIiHd3d2ZmZlVVVVVVVURERERERDMzM0RERDMzM0RERDMzMzMzMzMzMzMzMzMzM0RERERERCIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIiIiIjMzMyIiIhERESIiIhERESIiIiIiIjMzMzMzMzMzMyIiIjMzMzMzMyIiIiIiIhERERERESIiIiIiIjMzMzMzMyIiIhERESIiIhERESIiIiIiIjMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIhERESIiIiIiIjMzMzMzMyIiIjMzMzMzMyIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM0RERERERERERERERDMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMyIiIhERESIiIiIiIjMzMyIiIiIiIjMzMyIiIiIiIiIiIiIiIhERESIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIjMzMzMzMyIiIhERESIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIhERESIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIhERESIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERFVVVURERDMzMzMzM0RERERERERERDMzMzMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIhERERERERERESIiIhERERERESIiIiIiIiIiIiIiIiIiIhERESIiIhERERERESIiIhERESIiIiIiIhERESIiIhERESIiIhERESIiIhERERERESIiIhERESIiIiIiIkRERERERDMzM0RERERERDMzMzMzM0RERDMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIhERERERESIiIiIiIiIiIjMzMzMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIhERERERERERESIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIhERESIiIiIiIiIiIhERESIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIhERESIiIiIiIiIiIiIiIhERERERESIiIhERESIiIiIiIiIiIiIiIiIiIhERESIiIiIiIjMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERERERERERFVVVWZmZoiIiHd3d4iIiKqqqqqqqqqqqszMzO7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7u7u7////////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3MzMzMzMy7u7uqqqqqqqqqqqq7u7u7u7uqqqqZmZmZmZmZmZmqqqqqqqqqqqqqqqq7u7uqqqqqqqq7u7u7u7u7u7u7u7u7u7u7u7u7u7uZmZmIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3dVVVVmZmZmZmZmZmZVVVVmZmZmZmZVVVVVVVVVVVVERERVVVVERERVVVVERERERERVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZmqqqqZmZmqqqq7u7u7u7u7u7u7u7u7u7uqqqqZmZmZmZmZmZmZmZmZmZmZmZmZmZmIiIiIiIh3d3dmZmZmZmZmZmZmZmZVVVVmZmZVVVVVVVVVVVVmZmZ3d3dmZmZ3d3d3d3d3d3d3d3eIiIiZmZmqqqqZmZmqqqqZmZmZmZmZmZmZmZmZmZmqqqqZmZmIiIh3d3d3d3d3d3dmZmZmZmZmZmZ3d3d3d3dmZmZmZmZVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVmZmaZmZmIiIhmZmZVVVV3d3d3d3d3d3dmZmZVVVVEREQzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzNEREQzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMiIiIiIiIiIiIiIiIREREiIiIREREiIiIiIiIzMzMiIiIiIiIREREiIiIREREiIiIzMzMzMzMzMzMzMzMiIiIiIiIiIiIREREiIiIREREiIiIiIiJEREREREQiIiIREREREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIREREREREREREiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNEREQzMzMzMzNEREQzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIREREREREiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMiIiJEREQzMzMzMzMiIiIzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIiIiIREREiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIREREiIiIREREiIiIzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzNEREQzMzMzMzMzMzMzMzNEREREREQzMzNEREQzMzNEREREREREREQzMzMzMzNEREREREQzMzMiIiIzMzMiIiIzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIREREiIiIREREREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIREREiIiIREREiIiIREREREREiIiIiIiIREREREREiIiIiIiIREREiIiIiIiIREREiIiIiIiIzMzMzMzMzMzMzMzNERERVVVVEREQzMzNEREREREQzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIzMzMiIiIiIiIREREiIiIiIiIiIiIzMzMzMzMiIiIzMzMiIiIiIiIREREiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIREREiIiIREREiIiIiIiIREREiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzNERERERERVVVVVVVVmZmZ3d3eZmZmZmZmIiIiIiIiZmZm7u7vMzMzu7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u////////////7u7u7u7u////7u7u////7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3d7u7u3d3d7u7u3d3d3d3d3d3dzMzM3d3dzMzMu7u7u7u7qqqqmZmZiIiIiIiImZmZiIiIiIiId3d3d3d3ZmZmd3d3d3d3d3d3iIiImZmZmZmZqqqqqqqqqqqqqqqqqqqqqqqqu7u7u7u7qqqqmZmZqqqqqqqqqqqqqqqqmZmZqqqqiIiId3d3d3d3iIiId3d3ZmZmZmZmd3d3ZmZmVVVVREREVVVVREREVVVVREREREREVVVVREREVVVVVVVVVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmd3d3d3d3d3d3d3d3iIiIiIiId3d3iIiIiIiImZmZiIiIqqqqqqqqqqqqzMzMzMzMu7u7u7u7u7u7u7u7qqqqqqqqmZmZiIiIiIiIiIiId3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3iIiImZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZiIiIiIiId3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmZmZmVVVVVVVVREREVVVVREREVVVVVVVVREREVVVVVVVVREREREREREREREREREREREREZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmVVVVMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzIiIiMzMzERERERERERERIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiERERIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiERERERERIiIiERERMzMzMzMzIiIiIiIiERERERERIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzIiIiIiIiERERIiIiMzMzMzMzMzMzMzMzIiIiIiIiERERERERIiIiERERIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiERERERERIiIiIiIiIiIiIiIiERERIiIiMzMzIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREMzMzMzMzIiIiIiIiMzMzMzMzIiIiMzMzIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiERERERERERERIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiERERIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiMzMzMzMzMzMzIiIiMzMzMzMzIiIiMzMzMzMzMzMzIiIiIiIiERERERERIiIiMzMzMzMzIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREREREREREMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREREREREREREREREREMzMzMzMzIiIiMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiMzMzMzMzMzMzMzMzREREMzMzIiIiIiIiIiIiIiIiIiIiIiIiERERERERIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiERERERERIiIiIiIiERERIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzREREMzMzREREREREREREREREREREMzMzMzMzIiIiERERIiIiIiIiIiIiERERERERERERMzMzREREMzMzIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiERERIiIiERERIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzAP//AAAzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMiIiIzMzNEREQzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzNERERERERERERVVVVVVVVmZmaIiIiIiIiIiIiIiIiIiIiZmZm7u7vd3d3u7u7////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u7u7u////////////7u7u////////////7u7u7u7u7u7u////7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMu7u7u7u7u7u7u7u7u7u7qqqqmZmZmZmZiIiIiIiIiIiIZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmVVVVVVVVZmZmd3d3d3d3d3d3iIiImZmZiIiImZmZmZmZqqqqqqqqqqqqqqqqu7u7zMzMqqqqu7u7u7u7u7u7u7u7qqqqqqqqqqqqmZmZiIiIiIiImZmZiIiId3d3ZmZmZmZmVVVVREREVVVVREREVVVVREREVVVVVVVVREREVVVVREREREREREREREREREREREREREREREREREREREREVVVVVVVVREREREREVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3d3d3mZmZiIiImZmZqqqqmZmZmZmZqqqqqqqqu7u7u7u7zMzMzMzMu7u7u7u7qqqqqqqqmZmZiIiId3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3mZmZiIiImZmZiIiImZmZiIiImZmZiIiImZmZmZmZiIiIiIiIiIiId3d3ZmZmZmZmVVVVVVVVREREREREREREREREREREREREVVVVVVVVVVVVZmZmZmZmd3d3ZmZmVVVVVVVVVVVVREREVVVVVVVVVVVVREREREREREREREREMzMzREREMzMzREREREREREREMzMzVVVVZmZmVVVVVVVVREREREREIiIiMzMzMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiERERIiIiIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiERERIiIiERERERERIiIiIiIiMzMzIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiERERERERIiIiIiIiERERIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERERERIiIiERERERERERERMzMzMzMzIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiMzMzMzMzREREMzMzREREMzMzREREMzMzIiIiIiIiIiIiMzMzIiIiMzMzMzMzIiIiMzMzIiIiIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiERERIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiERERERERERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiMzMzIiIiMzMzMzMzIiIiMzMzIiIiIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiERERIiIiERERIiIiMzMzMzMzIiIiIiIiMzMzIiIiMzMzMzMzIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREMzMzIiIiMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiERERIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzREREREREREREREREREREREREMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERMzMzVVVVMzMzERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiERERERERERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiMzMzMzMzREREREREREREMzMzMzMzIiIiIiIiIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzREREREREIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREVVVVREREREREREREZmZmiIiId3d3d3d3d3d3d3d3d3d3mZmZu7u73d3d7u7u////////////////////////////7u7u////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////+7u7v///+7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7v///+7u7u7u7v///////+7u7v///+7u7v///+7u7v///////+7u7v///+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3czMzN3d3czMzMzMzLu7u7u7u6qqqqqqqqqqqpmZmZmZmXd3d3d3d3d3d3d3d3d3d1VVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d3d3d3d3d4iIiIiIiHd3d4iIiIiIiJmZmbu7u6qqqru7u7u7u7u7u8zMzLu7u6qqqru7u7u7u7u7u6qqqqqqqqqqqqqqqpmZmZmZmYiIiHd3d3d3d3d3d2ZmZmZmZmZmZnd3d2ZmZmZmZlVVVVVVVURERERERERERERERDMzM0RERERERERERERERERERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVXd3d3d3d4iIiIiIiJmZmZmZmYiIiJmZmaqqqqqqqqqqqru7u6qqqqqqqqqqqpmZmaqqqpmZmYiIiHd3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZnd3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVURERERERERERERERERERDMzM0RERFVVVVVVVWZmZlVVVWZmZmZmZlVVVVVVVVVVVURERERERFVVVURERERERERERDMzM0RERDMzMzMzM0RERDMzM0RERDMzM0RERERERERERERERDMzMyIiIjMzMyIiIjMzMzMzMyIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIjMzMyIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIhERESIiIiIiIhERESIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIhERESIiIiIiIiIiIhERESIiIjMzMyIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMyIiIhERERERESIiIhERESIiIiIiIiIiIhERERERESIiIhERESIiIiIiIjMzMzMzMyIiIjMzMzMzMyIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzM0RERDMzM0RERERERDMzMzMzMzMzMyIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIjMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzMyIiIjMzMzMzMyIiIhERESIiIiIiIjMzMzMzM0RERDMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMyIiIiIiIhERESIiIiIiIhERESIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMyIiIiIiIjMzMyIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMxERERERESIiIiIiIiIiIiIiIhERESIiIiIiIhERESIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMyIiIjMzM0RERERERDMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIkRERDMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIjMzMzMzMyIiIiIiIhERESIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzM0RERERERERERDMzM0RERFVVVURERDMzMyIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIlVVVVVVVTMzMyIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIhERERERERERERERERERESIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzM0RERDMzMyIiIjMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzM0RERERERDMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERGZmZmZmZnd3d2ZmZmZmZnd3d3d3d4iIiKqqqszMzN3d3e7u7u7u7v///////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////u7u7u7u7d3d3MzMy7u7u7u7vMzMzd3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7////u7u7////////u7u7////u7u7////u7u7////////u7u7////u7u7////u7u7u7u7u7u7u7u7d3d3d3d3d3d3MzMzd3d3MzMzMzMzMzMy7u7vMzMy7u7u7u7u7u7u7u7u7u7uZmZmIiIiIiIiIiIiIiIh3d3dVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3dmZmZmZmZ3d3eIiIiIiIiZmZmZmZmZmZmZmZmZmZmqqqqqqqq7u7u7u7vMzMy7u7uqqqqqqqq7u7u7u7uZmZmZmZmZmZmqqqqZmZmIiIiZmZmIiIiIiIiIiIiIiIiIiIh3d3dVVVVEREREREREREQzMzMzMzMzMzMzMzNEREQzMzNERERERERERERERERERERERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3d3d3eIiIiIiIiZmZmZmZmqqqqqqqqqqqqZmZmZmZmZmZmIiIiIiIh3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZ3d3d3d3eIiIh3d3d3d3d3d3eIiIh3d3eIiIh3d3eIiIh3d3d3d3d3d3d3d3dmZmZmZmZmZmZVVVVVVVVVVVVERERERERERERERERERERERERVVVVVVVVVVVVERERmZmZ3d3dmZmZVVVVVVVVVVVVEREREREQzMzMzMzMzMzNEREQzMzNEREQzMzMzMzNEREREREREREREREREREQzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMiIiIREREREREiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIREREiIiIiIiIiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIzMzNEREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzNEREREREREREREREQzMzMzMzMiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzNEREQzMzMzMzMiIiIiIiIiIiIzMzMiIiIREREiIiIiIiIiIiIzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMiIiIREREREREiIiIREREREREREREiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMiIiIiIiIzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMiIiIiIiIiIiIzMzMzMzMzMzNEREQzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIREREiIiIiIiIREREiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiJEREQzMzMiIiIzMzMzMzMiIiIiIiIiIiIREREREREiIiIiIiIiIiIzMzMzMzMzMzMiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMiIiIiIiIzMzMzMzMiIiIiIiIREREiIiIzMzMzMzMiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIREREiIiIiIiIREREiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREREREiIiIiIiIiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIREREiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzNEREQzMzMzMzMiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzNERERERERERERERERERERVVVVVVVVmZmZ3d3dmZmZ3d3d3d3eIiIiZmZmZmZm7u7vu7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u3d3d7u7u3d3d3d3dzMzMu7u7u7u7zMzM3d3dzMzMu7u7u7u7u7u7zMzM3d3d3d3d3d3d7u7u7u7u7u7u////7u7u////////////////////////7u7u////7u7u////7u7u7u7u3d3d7u7u3d3dzMzM3d3du7u7zMzMzMzMu7u7u7u7u7u7u7u7zMzMu7u7u7u7zMzMqqqqqqqqu7u7qqqqmZmZmZmZiIiId3d3ZmZmd3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiId3d3iIiId3d3iIiIiIiIiIiIiIiIiIiImZmZmZmZmZmZmZmZqqqqqqqqu7u7mZmZmZmZmZmZu7u7qqqqqqqqqqqqu7u7qqqqmZmZmZmZmZmZiIiId3d3ZmZmVVVVVVVVVVVVVVVVREREREREREREREREREREREREMzMzREREMzMzREREMzMzREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3d3d3iIiImZmZmZmZiIiIiIiIiIiIiIiId3d3d3d3ZmZmVVVVVVVVZmZmZmZmVVVVVVVVZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmd3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVREREREREREREVVVVREREREREREREREREREREZmZmZmZmVVVVd3d3iIiIZmZmREREMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREIiIiIiIiMzMzMzMzMzMzIiIiREREMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiERERERERIiIiIiIiIiIiERERIiIiIiIiERERIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzIiIiIiIiIiIiERERERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiMzMzMzMzREREMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREMzMzMzMzIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiIiIiMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzREREMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzIiIiMzMzMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiERERERERIiIiERERIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiERERMzMzMzMzIiIiMzMzIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiERERIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiMzMzREREIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzREREREREMzMzIiIiIiIiMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzIiIiIiIiREREREREREREMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiMzMzIiIiIiIiMzMzMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzIiIiMzMzMzMzIiIiMzMzMzMzMzMzMzMzIiIiIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzREREMzMzMzMzREREREREMzMzMzMzMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiERERIiIiIiIiERERIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiERERERERIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiERERIiIiERERERERIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzIiIiMzMzMzMzIiIiMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzREREREREREREVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3iIiIiIiIqqqq3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////+7u7u7u7u7u7v///+7u7v///////////+7u7u7u7u7u7t3d3czMzKqqqru7u8zMzN3d3d3d3d3d3d3d3e7u7u7u7u7u7u7u7v///+7u7u7u7v///+7u7v///+7u7v///+7u7v///+7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3bu7u7u7u7u7u7u7u7u7u7u7u8zMzMzMzMzMzLu7u7u7u7u7u7u7u6qqqqqqqru7u5mZmZmZmZmZmYiIiHd3d3d3d2ZmZnd3d2ZmZmZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZmZmZnd3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d2ZmZmZmZnd3d3d3d3d3d4iIiIiIiIiIiJmZmZmZmZmZmaqqqqqqqpmZmaqqqqqqqqqqqpmZmZmZmaqqqqqqqoiIiIiIiHd3d4iIiHd3d4iIiHd3d4iIiGZmZmZmZmZmZmZmZlVVVVVVVURERERERDMzM0RERDMzM0RERERERERERERERERERERERERERFVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d4iIiIiIiIiIiIiIiHd3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVWZmZnd3d4iIiIiIiJmZmZmZmZmZmYiIiHd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVURERFVVVURERFVVVURERFVVVVVVVURERFVVVURERERERERERFVVVURERERERFVVVWZmZoiIiHd3d1VVVTMzMyIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIjMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzM0RERDMzMyIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIiIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIjMzMyIiIhERESIiIhERESIiIiIiIjMzMyIiIiIiIiIiIjMzMyIiIiIiIjMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIiIiIiIiIkRERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIhERESIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERERERERERERERDMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMyIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzM0RERDMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIjMzMyIiIjMzMyIiIiIiIjMzMyIiIiIiIiIiIiIiIhERERERERERESIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIiIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzMyIiIjMzMzMzM1VVVURERDMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMyIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzM0RERERERFVVVURERDMzMzMzMyIiIjMzMzMzMzMzMyIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIjMzM0RERERERERERCIiIjMzMzMzMzMzMyIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzM0RERDMzMzMzMzMzMzMzM0RERERERDMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIiIiIjMzMyIiIjMzM0RERFVVVTMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIjMzMyIiIiIiIiIiIjMzMzMzM0RERDMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzM0RERERERERERERERDMzMzMzMzMzM0RERDMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzMyIiIhERESIiIhERERERERERERERESIiIjMzMzMzMyIiIiIiIiIiIhERERERESIiIhERERERESIiIhERESIiIhERERERESIiIhERESIiIiIiIiIiIhERESIiIiIiIiIiIiIiIhERERERESIiIhERERERESIiIhERESIiIhERESIiIiIiIiIiIjMzMyIiIjMzMzMzMyIiIiIiIiIiIhERESIiIhERESIiIhERERERESIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIiIiIjMzMyIiIjMzMzMzMyIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzM0RERERERFVVVVVVVURERERERFVVVVVVVWZmZmZmZmZmZmZmZnd3d5mZmbu7u8zMzN3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7d3d3d3d3d3d3d3d3d3d3MzMzMzMzd3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7////////////u7u7////u7u7u7u7////u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzd3d3MzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7uqqqqZmZmZmZmIiIiIiIiZmZmIiIiIiIiZmZmIiIh3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3eIiIiIiIiIiIiIiIiIiIiZmZmIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3eIiIiIiIiZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmIiIiIiIiIiIiIiIiIiIiZmZmZmZmIiIiIiIiIiIiIiIiIiIhmZmZmZmZVVVVVVVVVVVVERERERERERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZmZmZ3d3d3d3d3d3d3d3dmZmZmZmZmZmZVVVVmZmZVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVmZmZ3d3eIiIiZmZmqqqqZmZmZmZmZmZmIiIiIiIh3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVERERVVVVERERERERERERERERERERERERERERERERERERERERERERERERERERVVVVmZmZmZmZmZmZ3d3d3d3dmZmZEREQzMzMzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzNEREQzMzMzMzMzMzMzMzMiIiIiIiIiIiIzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIREREiIiIzMzMiIiIiIiIiIiIREREiIiIiIiIREREiIiIzMzMiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzNEREREREQzMzMzMzMzMzNEREQzMzMzMzMzMzMiIiIREREiIiIiIiIREREiIiIiIiIzMzMiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMREREzMzMzMzMzMzMiIiIiIiIzMzMiIiIzMzNEREQzMzNEREREREREREREREREREREREREREQzMzMiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIREREREREREREiIiIiIiIiIiIzMzMiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIzMzMzMzMzMzMiIiIREREiIiIiIiIzMzMiIiIzMzMiIiIiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzMzMzMzMzMiIiIiIiIzMzMiIiIiIiIzMzMiIiIzMzMiIiIiIiIzMzMiIiIzMzMzMzNEREQzMzMzMzMzMzNERERERERVVVUzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIzMzNVVVVVVVVEREQiIiIzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzNEREREREREREREREQzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzMiIiIiIiIzMzMiIiIiIiIiIiIzMzNEREQzMzMiIiIzMzMiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiJEREQzMzMiIiIiIiIiIiIzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNERERERERERERERERERERVVVVEREQzMzMzMzNEREQzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIiIiIREREREREiIiIREREiIiIREREREREzMzMiIiIiIiIREREREREiIiIREREREREiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIREREiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIREREiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzNEREQzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMzMzMiIiIzMzMiIiIzMzMiIiIiIiIzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzNERERERERERERERERERERERERVVVVVVVVmZmZVVVV3d3eIiIiZmZmqqqq7u7u7u7vd3d3u7u7////////////////u7u7////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////7u7u3d3dzMzMu7u7zMzMzMzMzMzMzMzM3d3d3d3d7u7u7u7u7u7u7u7u////7u7u////7u7u7u7u7u7u7u7u////7u7u7u7u////7u7u////7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMu7u7u7u7qqqqmZmZiIiIiIiIiIiIiIiImZmZmZmZiIiIiIiImZmZd3d3d3d3d3d3d3d3d3d3iIiId3d3iIiId3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3iIiIiIiId3d3ZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3iIiIiIiImZmZiIiIiIiImZmZqqqqqqqqmZmZqqqqqqqqqqqqiIiImZmZqqqqmZmZiIiIiIiIiIiIiIiId3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVd3d3d3d3iIiIiIiIiIiImZmZmZmZmZmZiIiIiIiId3d3ZmZmVVVVVVVVREREREREREREREREREREREREREREREREREREREREREREREREREREREREMzMzREREREREVVVVVVVVd3d3d3d3iIiId3d3ZmZmVVVVVVVVREREREREMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzREREREREVVVVREREMzMzMzMzIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiERERIiIiIiIiIiIiMzMzMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzREREMzMzMzMzIiIiMzMzREREMzMzMzMzERERERERIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiREREREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREMzMzREREREREREREREREREREREREMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiMzMzIiIiMzMzMzMzIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiIiIiIiIiERERERERIiIiIiIiIiIiIiIiERERIiIiERERERERIiIiERERIiIiIiIiIiIiREREREREREREMzMzMzMzIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzMzMzIiIiIiIiIiIiMzMzIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzREREVVVVMzMzMzMzMzMzREREREREMzMzIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiERERIiIiIiIiMzMzMzMzMzMzMzMzREREVVVVREREREREMzMzMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiMzMzREREIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzREREREREREREREREREREREREMzMzREREVVVVREREREREREREMzMzREREMzMzMzMzMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiERERERERIiIiERERERERIiIiIiIiIiIiERERIiIiERERERERIiIiERERERERIiIiIiIiIiIiERERIiIiIiIiERERIiIiIiIiIiIiMzMzIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiERERIiIiIiIiERERIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiMzMzMzMzMzMzIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzMzMzIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzREREREREREREREREREREZmZmZmZmZmZmd3d3iIiImZmZqqqqqqqqu7u73d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7t3d3bu7u7u7u7u7u8zMzN3d3d3d3d3d3e7u7u7u7u7u7v///+7u7u7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7v///+7u7u7u7v///////+7u7u7u7u7u7t3d3e7u7t3d3e7u7t3d3e7u7u7u7u7u7u7u7t3d3d3d3czMzN3d3czMzMzMzMzMzLu7u7u7u7u7u6qqqqqqqqqqqpmZmZmZmZmZmYiIiIiIiIiIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiJmZmZmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiIiIiHd3d2ZmZnd3d3d3d4iIiIiIiHd3d2ZmZlVVVVVVVVVVVURERERERERERFVVVURERERERERERERERERERFVVVVVVVVVVVWZmZnd3d4iIiIiIiJmZmaqqqqqqqru7u7u7u6qqqqqqqqqqqqqqqqqqqoiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVVVVVURERERERERERERERERERFVVVURERFVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVURERERERERERFVVVVVVVURERERERFVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZlVVVWZmZmZmZmZmZmZmZlVVVWZmZlVVVVVVVURERDMzMzMzMzMzM0RERDMzM0RERERERERERERERERERERERERERERERDMzMzMzM0RERDMzM0RERERERGZmZnd3d3d3d1VVVURERFVVVURERDMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERFVVVURERDMzMyIiIiIiIhERESIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIjMzMzMzMzMzMyIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzM0RERDMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM0RERERERERERERERFVVVTMzMyIiIiIiIiIiIjMzMyIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIhERESIiIhERERERESIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIkRERDMzMzMzMyIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMyIiIjMzMyIiIiIiIhERERERESIiIiIiIiIiIiIiIjMzMyIiIhERETMzM0RERDMzMzMzMzMzMyIiIjMzMyIiIiIiIhERERERESIiIiIiIiIiIiIiIhERERERERERESIiIiIiIiIiIhERESIiIiIiIjMzMyIiIiIiIkRERDMzMzMzMyIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIjMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIhERESIiIiIiIjMzMzMzM0RERCIiIiIiIjMzMzMzM0RERDMzMyIiIkRERDMzMyIiIiIiIiIiIhERESIiIhERESIiIhERERERERERESIiIiIiIjMzMzMzMzMzMzMzM0RERERERFVVVURERDMzMzMzMyIiIiIiIiIiIjMzMyIiIjMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMyIiIjMzM0RERERERCIiIiIiIiIiIjMzMyIiIiIiIhERESIiIiIiIiIiIhERERERESIiIjMzMyIiIiIiIjMzMyIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMyIiIiIiIhERETMzMzMzMzMzMzMzMzMzM0RERERERERERDMzM0RERERERERERERERERERERERDMzMzMzM0RERFVVVURERERERDMzMzMzMzMzMyIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIiIiIhERESIiIhERERERESIiIhERESIiIiIiIiIiIhERERERESIiIhERESIiIhERESIiIhERESIiIiIiIhERERERERERESIiIhERESIiIiIiIjMzMyIiIhERERERESIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIjMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIjMzM0RERDMzMyIiIiIiIiIiIhERERERESIiIiIiIiIiIiIiIjMzMzMzM0RERDMzM0RERERERERERFVVVVVVVVVVVWZmZmZmZnd3d3d3d5mZmaqqqru7u8zMzN3d3d3d3f///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3d3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7////////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7////u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3MzMzMzMy7u7uqqqqqqqqqqqqqqqqqqqqqqqqZmZmZmZmZmZmIiIiIiIiZmZmIiIiIiIiIiIiIiIh3d3d3d3eIiIiIiIiZmZmZmZmZmZmqqqqqqqq7u7uqqqqqqqqqqqqZmZmIiIiIiIiIiIiIiIiIiIh3d3d3d3dVVVVVVVVVVVVVVVVVVVVERERERERERERVVVVVVVVVVVVEREREREQzMzNERERERERERERVVVVmZmZmZmZ3d3d3d3eIiIiIiIiZmZmIiIiZmZmZmZmqqqqqqqqZmZmZmZmIiIiIiIiIiIh3d3d3d3d3d3eIiIh3d3d3d3dmZmZ3d3dmZmZmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVEREREREQzMzNEREQzMzNEREREREREREREREREREQzMzNERERVVVVERERERERVVVVERERERERERERERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVEREREREREREREREQzMzNEREQzMzNEREQzMzMzMzMzMzNEREREREREREREREREREREREREREQzMzMzMzMzMzMzMzNERERERERERERVVVVVVVVVVVVEREQzMzMzMzMiIiIiIiIzMzMiIiIzMzNEREREREQzMzNERERERERVVVUzMzMzMzMzMzNEREREREREREQzMzMiIiIiIiIREREiIiIzMzMiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMiIiIzMzMiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIzMzNEREQzMzMzMzMzMzMzMzMiIiJEREQzMzNEREQzMzMzMzMzMzNERERERERERERVVVVEREQzMzMiIiIzMzMiIiIzMzMiIiIREREREREiIiIREREREREiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMiIiIREREiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREREREREREQzMzMzMzNEREREREREREQiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIREREREREREREiIiIiIiIiIiIzMzMiIiIREREzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIzMzMiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiJERERVVVVEREQzMzMzMzMzMzMiIiIREREiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIzMzMzMzMzMzMiIiIiIiIREREiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIzMzMiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzMzMzMzMzNEREQzMzMzMzMiIiIzMzMiIiIiIiIzMzMiIiIzMzMiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIzMzMzMzNEREQzMzMiIiIiIiIzMzMzMzMzMzMzMzMiIiIiIiIREREiIiIiIiIiIiIREREREREiIiIREREiIiIiIiIiIiIiIiIzMzMzMzNEREREREQzMzNEREREREREREQzMzMzMzMiIiIzMzMzMzMiIiIzMzMzMzMiIiIzMzMiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzNEREREREQzMzMiIiIiIiIiIiIiIiIREREREREiIiIREREREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIzMzNEREREREQzMzMzMzMzMzMzMzNEREREREREREREREQzMzNEREQzMzNEREQzMzMzMzNVVVVmZmZmZmZVVVVEREQzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIREREREREiIiIREREREREiIiIREREiIiIiIiIREREiIiIREREREREiIiIREREiIiIREREiIiIREREREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzNEREREREQiIiIzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIzMzMiIiIiIiIzMzMiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIzMzMzMzNERERERERERERVVVVERERVVVVERERVVVVmZmZmZmZmZmZmZmaIiIiqqqq7u7uqqqq7u7vMzMzu7u7u7u7////////////////////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7uzMzM3d3d3d3d7u7u7u7u7u7u7u7u////////////////////////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u////////7u7u7u7u7u7u3d3d7u7u3d3dzMzMzMzMu7u7qqqqqqqqiIiIiIiImZmZmZmZiIiId3d3iIiIiIiImZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZmZmZiIiIiIiImZmZmZmZmZmZmZmZqqqqqqqqu7u7u7u7qqqqqqqqmZmZiIiIiIiId3d3ZmZmZmZmVVVVREREREREREREREREVVVVVVVVZmZmd3d3VVVVREREREREMzMzREREREREREREVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmd3d3d3d3iIiIiIiIiIiImZmZiIiIiIiId3d3iIiIiIiIiIiIiIiIZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREREREMzMzMzMzREREREREREREMzMzMzMzMzMzREREVVVVREREREREREREREREREREREREREREVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVREREREREREREREREREREMzMzREREREREREREMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVREREVVVVREREMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzREREVVVVVVVVREREVVVVREREMzMzREREMzMzMzMzMzMzIiIiERERERERIiIiMzMzMzMzIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzIiIiREREREREMzMzMzMzIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiMzMzIiIiMzMzREREMzMzMzMzMzMzIiIiIiIiIiIiERERMzMzMzMzMzMzREREMzMzIiIiMzMzMzMzMzMzREREMzMzMzMzREREMzMzREREREREMzMzREREMzMzMzMzIiIiIiIiIiIiIiIiERERERERERERIiIiIiIiERERIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiERERIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzREREREREREREVVVVREREREREREREREREMzMzMzMzREREREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREMzMzMzMzIiIiIiIiMzMzIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiREREMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzIiIiIiIiERERIiIiERERIiIiIiIiMzMzIiIiIiIiERERIiIiMzMzREREVVVVVVVVREREIiIiIiIiERERERERERERERERERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiMzMzMzMzREREMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzMzMzIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVREREREREMzMzREREREREMzMzMzMzMzMzIiIiIiIiIiIiMzMzIiIiIiIiMzMzIiIiIiIiMzMzMzMzIiIiMzMzIiIiMzMzREREMzMzIiIiIiIiIiIiMzMzMzMzREREMzMzMzMzIiIiERERERERIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzREREREREVVVVREREMzMzREREREREMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzIiIiERERERERIiIiERERERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzMzMzMzMzREREMzMzMzMzMzMzREREMzMzREREREREREREREREMzMzREREMzMzREREMzMzREREVVVVd3d3ZmZmREREMzMzMzMzMzMzREREREREMzMzMzMzIiIiIiIiIiIiIiIiERERERERIiIiERERIiIiERERIiIiIiIiERERIiIiERERERERIiIiERERERERERERIiIiIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiMzMzERERERERIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiIiIiIiIiIiIiMzMzMzMzREREREREREREMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiMzMzIiIiIiIiMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzMzMzREREVVVVREREVVVVREREREREREREVVVVVVVVZmZmZmZmZmZmd3d3mZmZmZmZqqqqqqqqzMzM7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7t3d3d3d3d3d3e7u7u7u7u7u7u7u7v///+7u7v///+7u7v///////////////////////+7u7u7u7v///+7u7v///+7u7u7u7u7u7u7u7t3d3d3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3czMzLu7u7u7u5mZmYiIiIiIiHd3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiIiIiHd3d3d3d2ZmZnd3d4iIiIiIiIiIiIiIiJmZmaqqqpmZmaqqqqqqqqqqqpmZmYiIiIiIiHd3d3d3d2ZmZnd3d2ZmZmZmZlVVVVVVVVVVVWZmZnd3d1VVVVVVVURERERERERERERERERERERERFVVVVVVVWZmZlVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d2ZmZnd3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d3d3d2ZmZmZmZlVVVURERERERFVVVVVVVURERFVVVURERERERERERERERERERERERFVVVURERERERFVVVVVVVURERERERERERFVVVVVVVWZmZmZmZlVVVWZmZlVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVVVVVXd3d2ZmZkRERERERDMzMzMzMzMzM0RERDMzMyIiIjMzMzMzMzMzM0RERERERERERFVVVVVVVTMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMzMzM0RERDMzM0RERERERERERERERERERDMzMzMzMzMzMyIiIjMzMyIiIiIiIhERETMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIjMzMzMzMzMzMyIiIiIiIjMzM0RERGZmZlVVVTMzMyIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIkRERDMzMzMzMyIiIjMzMzMzM0RERDMzM0RERDMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIhERESIiIhERESIiIiIiIjMzMzMzMzMzM0RERDMzM0RERERERERERERERFVVVTMzMzMzMzMzMzMzM0RERDMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIjMzMyIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzM0RERFVVVURERDMzMzMzMyIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzM1VVVURERCIiIiIiIhERESIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMzMzMzMzMzMzM0RERERERERERDMzMzMzMzMzMzMzMzMzM0RERERERDMzMyIiIjMzMzMzMyIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVVVVVURERDMzM0RERERERFVVVVVVVTMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMyIiIjMzMzMzMyIiIjMzMyIiIjMzM0RERERERDMzMzMzMzMzMzMzMyIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIkRERERERERERERERERERERERERERERERDMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVURERDMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIhERESIiIhERERERESIiIiIiIiIiIhERESIiIhERERERERERESIiIhERESIiIhERESIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERDMzMzMzM0RERERERERERCIiIjMzM2ZmZnd3d1VVVURERERERERERERERDMzMzMzMzMzMyIiIiIiIiIiIhERERERESIiIhERESIiIhERERERERERESIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIhERERERESIiIiIiIhERERERESIiIhERERERETMzMyIiIiIiIiIiIiIiIhERESIiIhERERERESIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIjMzM0RERDMzMzMzMzMzMzMzMyIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMyIiIiIiIiIiIjMzMzMzMyIiIjMzMyIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIhERESIiIiIiIjMzMzMzMyIiIhERESIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzM0RERERERERERDMzMzMzM0RERFVVVURERFVVVVVVVWZmZmZmZnd3d4iIiJmZmaqqqru7u8zMzN3d3e7u7v///////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////u7u7d3d3MzMzMzMzd3d3d3d3u7u7u7u7u7u7////////////////u7u7////////u7u7////////////////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7d3d3d3d3MzMzMzMy7u7uqqqqIiIh3d3dmZmZVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVERERVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZmZmZ3d3eIiIh3d3d3d3eIiIiIiIh3d3eZmZmIiIiIiIiIiIiIiIh3d3eIiIiIiIiIiIiIiIh3d3dmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERERERERERERERVVVVERERmZmZmZmZ3d3dVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVERERERERERERERERERERERERmZmZVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVWIiIiIiIh3d3dmZmZEREREREREREREREREREQzMzMzMzMzMzNEREQzMzNEREQzMzNEREREREQzMzMzMzMzMzMiIiIiIiIzMzMiIiIzMzMzMzMiIiIzMzNEREQzMzMzMzNEREQzMzMzMzMiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVVVVVEREQzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREQzMzMzMzMzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIREREzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERVVVVEREQzMzMzMzMzMzNEREREREQzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIzMzMzMzMiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIzMzMzMzMiIiIzMzMiIiIiIiIiIiIzMzMzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIzMzMzMzNmZmZmZmZEREQzMzMiIiIiIiIzMzMiIiIiIiIiIiIzMzMiIiIzMzMiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIzMzMiIiIzMzMiIiIzMzMzMzMzMzNEREQzMzNEREREREQzMzMzMzMzMzMzMzNERERERERVVVVmZmZEREQzMzMiIiIzMzMzMzMzMzMzMzMzMzNEREQzMzNERERERERERERERERVVVVmZmZVVVVEREREREQzMzNERERERERVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzMzMzMzMzMzMzMiIiIiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzNERERERERVVVVVVVVEREREREQzMzMzMzNEREQzMzNEREREREREREREREREREREREQzMzMzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIREREiIiIREREREREREREREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIzMzMiIiIiIiIzMzMiIiIiIiIzMzMzMzMiIiIzMzMzMzNEREREREREREREREQzMzMzMzNERERVVVVVVVVEREQzMzMzMzNVVVVmZmZmZmZVVVVEREREREQzMzMzMzMiIiIiIiIiIiIREREREREiIiIREREiIiIREREREREiIiIREREiIiIiIiIiIiIiIiIREREREREiIiIREREiIiIREREiIiIiIiIiIiIREREiIiIiIiIiIiIREREiIiIiIiIzMzMiIiIREREREREiIiIREREiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzMiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIREREREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzNEREREREQzMzMzMzNERERERERERERERERVVVVmZmZVVVVmZmZ3d3d3d3eIiIiZmZmqqqq7u7vd3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3d3d3dzMzMzMzM3d3d3d3d7u7u7u7u7u7u7u7u7u7u////////////////////////7u7u////7u7u////7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u7u7u3d3d7u7u7u7u7u7u3d3dzMzMqqqqqqqqmZmZiIiIZmZmVVVVVVVVVVVVREREVVVVVVVVVVVVREREREREMzMzREREVVVVREREREREVVVVVVVVVVVVZmZmZmZmd3d3ZmZmiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3iIiIiIiIiIiIiIiImZmZiIiIiIiIiIiIiIiId3d3ZmZmZmZmVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmd3d3ZmZmVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3ZmZmZmZmZmZmVVVVREREVVVVVVVVREREVVVVREREREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVREREVVVVVVVVREREVVVVVVVVREREVVVVVVVVZmZmZmZmZmZmmZmZd3d3ZmZmVVVVVVVVVVVVREREMzMzMzMzIiIiMzMzMzMzREREMzMzMzMzMzMzREREMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiMzMzIiIiIiIiIiIiERERMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREREREMzMzREREREREREREMzMzREREMzMzMzMzMzMzMzMzREREREREREREREREREREREREVVVVREREREREMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREIiIiERERIiIiIiIiMzMzMzMzIiIiIiIiERERIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzMzMzREREMzMzMzMzMzMzREREREREREREREREREREREREMzMzMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzIiIiIiIiMzMzREREMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzIiIiIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzVVVVREREMzMzIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiERERIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzIiIiMzMzVVVVVVVVMzMzMzMzIiIiIiIiIiIiMzMzMzMzIiIiMzMzMzMzREREREREREREVVVVVVVVVVVVREREREREREREREREREREREREVVVVZmZmVVVVMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVREREREREVVVVREREVVVVREREREREMzMzMzMzMzMzIiIiMzMzREREREREREREREREREREVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREREREMzMzMzMzREREVVVVREREVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVREREREREMzMzREREMzMzREREREREVVVVREREVVVVREREREREREREREREREREVVVVREREREREREREREREREREREREREREREREREREREREMzMzMzMzMzMzREREMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiMzMzIiIiMzMzMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzIiIiIiIiMzMzREREREREMzMzMzMzREREREREREREREREMzMzREREREREVVVVREREMzMzREREZmZmiIiIZmZmVVVVREREREREMzMzIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERERERIiIiERERERERIiIiMzMzIiIiERERIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzREREREREREREREREREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiERERIiIiIiIiIiIiIiIiMzMzMzMzIiIiERERIiIiERERIiIiIiIiIiIiIiIiERERIiIiIiIiMzMzIiIiIiIiMzMzMzMzMzMzMzMzMzMzREREREREREREREREVVVVZmZmZmZmd3d3d3d3d3d3mZmZmZmZqqqqzMzM7u7u////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////+7u7u7u7u7u7t3d3d3d3d3d3d3d3e7u7u7u7u7u7v///////////////////////////////+7u7v///////+7u7v///+7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7t3d3e7u7t3d3e7u7t3d3e7u7u7u7u7u7u7u7t3d3d3d3d3d3bu7u7u7u6qqqoiIiIiIiGZmZlVVVURERERERFVVVVVVVURERERERERERERERERERERERFVVVVVVVWZmZmZmZnd3d3d3d4iIiIiIiIiIiHd3d4iIiIiIiIiIiIiIiIiIiHd3d4iIiHd3d3d3d2ZmZoiIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiGZmZnd3d3d3d2ZmZmZmZmZmZlVVVVVVVXd3d4iIiGZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZlVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZlVVVURERFVVVURERERERERERERERERERERERERERFVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVVVVVVVVVURERERERDMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERFVVVURERFVVVURERFVVVURERFVVVURERFVVVURERGZmZoiIiGZmZnd3d4iIiJmZmYiIiFVVVURERFVVVURERDMzMyIiIjMzMyIiIiIiIjMzMzMzMzMzMzMzM1VVVURERDMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzM0RERDMzMyIiIjMzM0RERDMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERERERERERDMzM0RERERERERERDMzM0RERERERERERDMzMzMzM0RERERERERERERERERERFVVVVVVVVVVVURERERERERERERERDMzMzMzMzMzM0RERDMzM0RERDMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERDMzMzMzM0RERERERDMzMyIiIiIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIjMzMzMzMzMzM0RERDMzM0RERDMzMzMzM0RERERERERERERERERERDMzMzMzM0RERERERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMyIiIjMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIkRERERERDMzM0RERERERDMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIiIiIjMzMyIiIiIiIjMzMzMzMzMzMzMzM0RERDMzMyIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMyIiIhERESIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzM0RERFVVVVVVVVVVVURERDMzM0RERDMzM0RERFVVVVVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERFVVVVVVVVVVVWZmZlVVVVVVVURERERERERERDMzM0RERFVVVWZmZkRERDMzMzMzM0RERDMzM0RERERERERERFVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVURERERERERERDMzM1VVVWZmZnd3d1VVVURERDMzMzMzMzMzMzMzM0RERFVVVVVVVURERFVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZlVVVVVVVURERERERERERGZmZnd3d1VVVVVVVTMzM0RERDMzMzMzMzMzMzMzM0RERFVVVVVVVWZmZnd3d3d3d2ZmZlVVVURERFVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVVVVVVVVVVVVVURERERERERERERERERERFVVVVVVVURERERERDMzMzMzMzMzM0RERERERERERERERDMzMzMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIiIiIjMzMzMzMzMzMyIiIjMzM0RERFVVVTMzM0RERERERERERERERDMzM0RERERERERERERERERERFVVVURERHd3d4iIiGZmZjMzMzMzMzMzMzMzMyIiIjMzMyIiIhERESIiIhERERERESIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIhERETMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIhERESIiIjMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzM0RERDMzMzMzMyIiIiIiIiIiIiIiIjMzM0RERCIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIhERESIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMyIiIhERERERESIiIiIiIiIiIiIiIjMzMyIiIiIiIhERESIiIhERESIiIhERERERESIiIiIiIiIiIhERERERESIiIiIiIjMzMzMzMzMzMyIiIjMzMzMzM0RERERERERERFVVVURERFVVVWZmZmZmZmZmZmZmZmZmZnd3d5mZmaqqqru7u8zMzO7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7d3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7////u7u7////////u7u7////////u7u7////////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMy7u7u7u7uZmZmIiIh3d3dmZmZERERERERERERVVVUzMzNERERERERERERVVVVVVVVmZmZ3d3eIiIiZmZmZmZmIiIiZmZmIiIh3d3eIiIh3d3eIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3dmZmZmZmZmZmZmZmZ3d3dmZmZmZmZ3d3d3d3eIiIiIiIh3d3d3d3eIiIiZmZmIiIiIiIh3d3d3d3d3d3dmZmZ3d3dmZmZmZmZmZmZ3d3d3d3dmZmZmZmZVVVVVVVVERERERERVVVVERERVVVVERERERERERERVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVERERERERERERERERVVVVVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZ3d3d3d3dmZmZmZmZVVVVVVVVEREREREQzMzNEREQzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzNEREQzMzNERERERERERERERERERERERERERERERERERERVVVV3d3eIiIh3d3eIiIiZmZmZmZlVVVVEREREREREREQzMzMzMzMzMzNEREQzMzNEREQzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIzMzNERERVVVVVVVVEREQzMzMzMzMzMzNEREQzMzMzMzNEREREREREREREREQzMzNEREREREREREQzMzMzMzMzMzNEREREREQzMzNERERERERERERERERERERERERVVVVmZmZVVVVVVVVEREREREREREREREREREREREREREREREQzMzMiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzNEREREREREREQzMzNEREQzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIiIiIzMzMiIiIzMzMiIiIiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIREREiIiIiIiIzMzNEREQzMzNEREQzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzNERERVVVUzMzNEREREREREREQzMzMiIiIiIiIzMzMzMzNVVVVEREQzMzNEREREREREREREREQzMzMiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIREREiIiIiIiIzMzNmZmZmZmZEREQzMzMiIiIiIiIiIiIREREiIiIREREiIiIiIiIzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIiIiIzMzNERERmZmZmZmZVVVUzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMiIiIzMzNEREQzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMiIiIiIiIzMzMzMzMiIiIzMzNERERERERVVVVVVVVmZmZ3d3dmZmZVVVVVVVVEREREREQzMzNERER3d3dmZmZVVVVEREQzMzMzMzMzMzMzMzMzMzNERERERERERERERERERERVVVVVVVVVVVVERERERERERERERERERERERERVVVVVVVVmZmZVVVVERERVVVVERERERERERERERERERERERERERERERERERERERERVVVVVVVUzMzNERERERERERERVVVVERERERERmZmZ3d3dmZmZVVVUzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVERERVVVVERERVVVVVVVVERERVVVVERERmZmZ3d3dmZmZEREREREREREREREREREQzMzNERERERERVVVVmZmZmZmZ3d3eIiIhmZmZVVVVmZmZVVVVmZmZVVVVVVVVVVVVmZmZ3d3dmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVERERERERERERERERVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIzMzMiIiIiIiJEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzNEREQzMzMzMzMzMzNERERERERERERERERVVVVERERVVVVERERERERVVVVVVVVmZmZVVVVEREQiIiIiIiIiIiIzMzMiIiIzMzMiIiIiIiIREREiIiIREREREREiIiIREREREREiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMiIiIREREiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIREREREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzNERERERERVVVVVVVVVVVVVVVVVVVVERERERERERERVVVVmZmZ3d3eIiIiZmZmZmZm7u7vMzMzu7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u////7u7u////////7u7u////////7u7u////////7u7u////7u7u7u7u////7u7u7u7u7u7u7u7u7u7u3d3d7u7u7u7u3d3d7u7u3d3d7u7u3d3d3d3d3d3dzMzMzMzMu7u7zMzMu7u7u7u7qqqqqqqqmZmZd3d3ZmZmVVVVVVVVREREREREREREVVVVREREVVVVVVVVVVVVd3d3iIiIqqqqmZmZmZmZiIiIiIiId3d3iIiIiIiId3d3iIiId3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmd3d3ZmZmZmZmVVVVZmZmZmZmZmZmd3d3d3d3d3d3mZmZmZmZmZmZmZmZmZmZmZmZmZmZqqqqmZmZmZmZmZmZd3d3iIiIiIiIZmZmZmZmZmZmVVVVVVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREREREREREVVVVVVVVREREREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVREREREREREREREREREREREREMzMzMzMzMzMzREREREREMzMzMzMzMzMzREREMzMzREREREREREREREREVVVVREREREREVVVVVVVVVVVVZmZmd3d3iIiIiIiIiIiIVVVVREREMzMzREREMzMzMzMzMzMzMzMzREREREREMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzMzMzREREREREREREREREMzMzMzMzMzMzREREREREREREREREREREREREREREREREREREMzMzMzMzMzMzREREMzMzREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVREREREREVVVVREREVVVVZmZmVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREMzMzMzMzIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzREREMzMzMzMzMzMzREREMzMzMzMzMzMzIiIiIiIiMzMzMzMzREREREREVVVVREREREREREREREREREREMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiERERERERIiIiIiIiIiIiREREVVVVMzMzIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzREREVVVVREREREREMzMzMzMzIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREREREVVVVREREMzMzMzMzMzMzIiIiMzMzMzMzREREMzMzREREREREMzMzMzMzREREREREREREREREREREMzMzREREREREMzMzREREZmZmZmZmREREMzMzMzMzIiIiIiIiIiIiMzMzVVVVREREMzMzREREREREREREREREREREREREREREREREMzMzMzMzREREMzMzREREVVVVREREREREREREREREREREREREREREREREMzMzMzMzREREREREREREREREREREMzMzREREMzMzREREVVVVMzMzMzMzREREVVVVREREREREMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzVVVVZmZmVVVVREREREREMzMzREREREREMzMzREREREREREREREREREREREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREd3d3iIiIZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3d3d3VVVVVVVVREREREREVVVVVVVVVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVREREMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzREREMzMzREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiERERIiIiIiIiMzMzMzMzMzMzIiIiIiIiERERIiIiIiIiERERIiIiIiIiIiIiMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiERERERERIiIiERERIiIiERERERERIiIiERERIiIiMzMzIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzREREREREREREREREREREREREREREREREVVVVZmZmd3d3iIiIiIiIiIiIiIiImZmZzMzM7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////+7u7v///////////////////////+7u7v///////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7v///+7u7v///////////+7u7v///+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3d3d3d3d3d3d3czMzMzMzMzMzLu7u7u7u7u7u5mZmYiIiIiIiHd3d2ZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVWZmZmZmZoiIiIiIiJmZmYiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d2ZmZmZmZlVVVWZmZlVVVURERFVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZnd3d3d3d4iIiIiIiIiIiIiIiJmZmYiIiJmZmaqqqqqqqru7u7u7u6qqqpmZmYiIiIiIiHd3d2ZmZmZmZlVVVVVVVVVVVURERFVVVVVVVVVVVURERFVVVVVVVVVVVURERFVVVURERERERERERDMzM0RERERERERERERERERERERERERERFVVVWZmZmZmZnd3d2ZmZmZmZlVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERDMzMzMzMzMzMzMzM0RERERERERERERERERERERERERERERERERERERERGZmZoiIiHd3d1VVVURERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzM0RERERERDMzMyIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIjMzM0RERDMzMzMzMzMzMzMzMzMzM0RERERERERERFVVVVVVVVVVVURERERERERERDMzMzMzMzMzM0RERERERERERERERERERERERERERFVVVVVVVVVVVVVVVURERFVVVURERFVVVWZmZmZmZnd3d2ZmZlVVVURERDMzMyIiIjMzMzMzMzMzMzMzM0RERERERERERERERDMzM0RERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMyIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIhERESIiIiIiIjMzMzMzMzMzMzMzMyIiIkRERDMzMzMzMzMzM0RERERERERERDMzM0RERDMzM0RERDMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERDMzM0RERDMzMzMzMzMzMyIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIhERESIiIjMzMyIiIjMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzMzMzM0RERDMzM0RERFVVVVVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIlVVVVVVVURERDMzMyIiIiIiIiIiIiIiIjMzM0RERERERDMzMzMzMzMzMzMzM0RERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzM1VVVURERERERDMzMzMzMzMzM0RERERERERERERERERERDMzM0RERERERDMzM0RERERERERERERERERERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIiIiIjMzMzMzM0RERFVVVURERERERDMzMzMzM0RERDMzM0RERDMzMzMzMzMzM0RERERERERERERERFVVVVVVVURERDMzM0RERERERERERERERFVVVWZmZmZmZlVVVURERFVVVVVVVVVVVWZmZlVVVVVVVWZmZlVVVWZmZmZmZnd3d3d3d2ZmZlVVVVVVVURERFVVVWZmZmZmZlVVVVVVVTMzM0RERDMzMzMzM0RERERERDMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzM0RERFVVVURERERERDMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzM0RERDMzM0RERDMzM0RERERERERERERERFVVVURERFVVVVVVVVVVVVVVVVVVVURERERERDMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzM0RERDMzMzMzMyIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzM0RERERERERERERERERERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIhERERERESIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIhERERERESIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIhERESIiIjMzMyIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIhERERERERERESIiIhERERERESIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzM0RERERERFVVVTMzMzMzM0RERERERERERFVVVWZmZnd3d4iIiIiIiIiIiJmZmczMzO7u7u7u7v///+7u7v///////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////u7u7////////////////////////u7u7////////////u7u7////////////////////////u7u7////////////////u7u7////////////////////u7u7////////////////////////////////////////////u7u7////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////u7u7////u7u7u7u7u7u7d3d3u7u7d3d3u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3MzMzMzMzMzMy7u7uqqqqqqqqZmZmIiIh3d3eIiIiIiIhmZmZ3d3eIiIh3d3dmZmZ3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVERERERERVVVVVVVVERERERERVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVV3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3dmZmZ3d3d3d3dmZmZVVVVVVVVVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERVVVVmZmZmZmZ3d3d3d3d3d3dmZmZVVVVmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVERERVVVVERERVVVVERERVVVVVVVVVVVVVVVVEREREREREREREREQzMzNERERERERVVVVVVVVVVVVVVVVEREREREQzMzMzMzMzMzNEREREREQzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzNERERERERERERVVVVmZmZVVVUzMzMzMzMzMzMzMzMiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIzMzMzMzMzMzMiIiIzMzMzMzNEREQzMzNERERERERERERVVVVVVVVmZmZmZmZVVVVEREQzMzMzMzNERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3eIiIhmZmZVVVVEREQzMzMzMzMzMzNEREREREREREREREREREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzNEREREREQzMzNEREREREREREQzMzMzMzMzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzNEREQzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMiIiIiIiIiIiIzMzMiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzNERERERERERERERERERERERERVVVVVVVVEREREREREREREREQzMzNEREQzMzMzMzNERERERERVVVVVVVVVVVVmZmZmZmZmZmZmZmZEREREREQzMzMzMzMzMzMzMzNVVVVVVVVEREQzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIzMzMzMzNEREREREREREQzMzMiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREREREQzMzMzMzNEREQzMzNEREREREREREREREQzMzMzMzNERERERERVVVVEREQzMzNEREREREREREREREQzMzNEREREREQzMzMzMzNEREREREQzMzNEREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIzMzMiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIzMzMzMzMzMzNEREREREREREREREREREREREREREREREREREREREQzMzNEREQzMzNERERERERERERERERVVVVVVVVEREREREREREREREREREQzMzNERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3dmZmZmZmZERERERERERERERERVVVVERERVVVVVVVVVVVVERERVVVVVVVVEREREREQzMzNERERERERVVVVVVVUzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREREREQzMzNERERERERERERERERVVVVVVVVERERVVVVVVVVEREREREREREREREQzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiJERERVVVVVVVVEREQzMzMzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzNEREREREREREREREREREQzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzNEREREREQzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIREREiIiIzMzMiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIREREiIiIiIiIiIiIREREREREiIiIiIiIREREiIiIREREiIiIREREiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzNEREQzMzMzMzMzMzNVVVVVVVVERERVVVVVVVVmZmaIiIiZmZmIiIiZmZmqqqrMzMzd3d3u7u7u7u7////////////////////////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u7u7u7u7u7u7u7u7u3d3d3d3dzMzM3d3d3d3d3d3d7u7u3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3dzMzMzMzMu7u7u7u7u7u7qqqqiIiIiIiImZmZd3d3iIiImZmZmZmZd3d3mZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmVVVVREREVVVVREREREREREREVVVVVVVVREREREREREREREREREREREREMzMzREREMzMzREREREREREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmVVVVZmZmd3d3d3d3iIiIiIiIiIiImZmZmZmZqqqqmZmZiIiImZmZmZmZmZmZmZmZiIiId3d3d3d3ZmZmVVVVVVVVVVVVVVVVREREREREREREREREMzMzREREREREREREVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVZmZmiIiId3d3VVVVREREVVVVREREREREREREREREREREREREVVVVREREREREREREIiIiMzMzMzMzMzMzREREREREREREIiIiMzMzIiIiMzMzMzMzMzMzMzMzREREMzMzMzMzREREVVVVZmZmVVVVVVVVMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzREREIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiMzMzREREREREMzMzREREREREVVVVREREVVVVZmZmZmZmVVVVVVVVREREMzMzMzMzREREREREREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmZmZmd3d3ZmZmZmZmd3d3d3d3ZmZmVVVVREREMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzIiIiMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzREREMzMzMzMzREREVVVVMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzMzMzREREMzMzMzMzIiIiIiIiIiIiERERIiIiMzMzIiIiERERIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzVVVVREREREREVVVVREREREREVVVVd3d3VVVVREREREREREREMzMzREREREREREREVVVVVVVVVVVVVVVVVVVVZmZmd3d3ZmZmZmZmVVVVREREREREREREMzMzIiIiREREVVVVREREMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiMzMzMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzVVVVREREREREREREREREMzMzREREREREREREREREREREMzMzREREMzMzREREREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzREREREREREREMzMzMzMzMzMzREREMzMzIiIiMzMzMzMzMzMzIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzMzMzREREREREREREREREREREREREREREREREMzMzMzMzREREMzMzREREREREREREREREVVVVREREREREREREREREREREMzMzREREREREREREVVVVREREREREREREREREVVVVVVVVREREVVVVREREVVVVREREVVVVZmZmVVVVZmZmVVVVVVVVREREVVVVVVVVZmZmVVVVZmZmd3d3ZmZmVVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmREREREREREREREREVVVVVVVVVVVVREREREREREREREREMzMzREREREREMzMzREREREREREREVVVVREREREREREREREREREREREREREREVVVVREREVVVVREREREREMzMzMzMzMzMzREREREREMzMzMzMzMzMzIiIiMzMzIiIiIiIiMzMzIiIiIiIiIiIiMzMzIiIiMzMzREREVVVVREREMzMzMzMzIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzREREMzMzREREREREMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzREREMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiERERERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzIiIiIiIiERERIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiERERERERIiIiIiIiERERERERIiIiIiIiIiIiERERERERIiIiERERIiIiERERERERIiIiIiIiERERERERERERERERIiIiERERERERIiIiIiIiIiIiMzMzMzMzMzMzREREMzMzIiIiMzMzMzMzVVVVVVVVREREVVVVVVVVZmZmd3d3iIiIiIiIiIiImZmZu7u7u7u73d3d7u7u7u7u////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7u7u7t3d3d3d3d3d3d3d3czMzN3d3czMzMzMzN3d3d3d3e7u7t3d3e7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3czMzLu7u7u7u7u7u6qqqpmZmaqqqoiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiJmZmZmZmZmZmZmZmZmZmYiIiIiIiIiIiHd3d3d3d2ZmZmZmZlVVVVVVVVVVVURERERERERERERERERERERERDMzM0RERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERERERFVVVVVVVWZmZlVVVVVVVWZmZmZmZmZmZmZmZnd3d4iIiJmZmZmZmaqqqpmZmZmZmZmZmZmZmZmZmaqqqpmZmYiIiIiIiHd3d3d3d2ZmZmZmZmZmZmZmZlVVVWZmZmZmZlVVVURERERERFVVVVVVVVVVVVVVVVVVVURERERERERERFVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZlVVVVVVVVVVVURERFVVVWZmZlVVVVVVVWZmZoiIiIiIiHd3d2ZmZlVVVVVVVURERDMzMzMzM0RERERERERERERERERERERERDMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzM0RERFVVVURERERERDMzM0RERFVVVVVVVVVVVURERDMzMyIiIiIiIjMzMzMzMyIiIjMzMyIiIjMzM0RERDMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIjMzM0RERDMzM0RERERERFVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZlVVVURERDMzM0RERERERERERERERERERFVVVWZmZmZmZmZmZmZmZlVVVWZmZnd3d2ZmZlVVVURERFVVVVVVVVVVVVVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzM0RERDMzMzMzM1VVVVVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIkRERDMzM0RERCIiIiIiIiIiIiIiIjMzMyIiIhERESIiIiIiIhERESIiIiIiIhERESIiIiIiIhERESIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVWZmZmZmZlVVVURERDMzM0RERGZmZmZmZmZmZlVVVURERERERERERFVVVURERFVVVVVVVVVVVVVVVURERERERFVVVVVVVVVVVTMzMzMzMzMzMzMzMzMzMyIiIjMzM0RERDMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIhERESIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERDMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERDMzM0RERFVVVURERERERDMzMzMzMzMzM0RERDMzMzMzM0RERERERERERDMzM0RERDMzM0RERDMzMzMzMzMzM0RERERERERERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzM0RERFVVVURERERERERERERERERERERERERERERERDMzM0RERERERERERERERERERERERERERERERERERERERERERDMzM0RERERERERERFVVVURERERERERERFVVVVVVVVVVVURERFVVVURERFVVVURERFVVVVVVVVVVVWZmZlVVVVVVVURERERERERERERERERERERERGZmZnd3d1VVVVVVVURERERERERERFVVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d3d3d2ZmZmZmZkRERERERFVVVVVVVVVVVURERERERERERERERERERERERERERERERERERERERFVVVVVVVURERERERFVVVVVVVURERERERFVVVVVVVURERERERERERERERDMzMzMzMzMzM0RERDMzM0RERDMzMzMzMzMzMyIiIiIiIjMzMzMzMyIiIiIiIjMzMyIiIjMzMzMzM0RERFVVVURERDMzMzMzMyIiIjMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM0RERDMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIjMzMzMzMyIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIhERESIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMyIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIhERERERESIiIhERESIiIiIiIiIiIhERESIiIhERESIiIhERESIiIhERESIiIhERESIiIiIiIiIiIjMzMzMzMzMzM0RERCIiIiIiIjMzM0RERERERERERERERERERFVVVVVVVWZmZnd3d3d3d4iIiJmZmaqqqru7u7u7u93d3f///+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7d3d3d3d3MzMy7u7u7u7vMzMzd3d3u7u7u7u7u7u7d3d3u7u7u7u7u7u7d3d3u7u7d3d3MzMzMzMy7u7uqqqqqqqq7u7uZmZmIiIiZmZmZmZmIiIiIiIiZmZl3d3d3d3d3d3eIiIh3d3eIiIiIiIiIiIiqqqqqqqqZmZmZmZmIiIiIiIh3d3d3d3dmZmZVVVVVVVVERERVVVVEREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzNERERERERERERERERERERERERVVVVmZmZVVVVmZmZVVVV3d3eIiIiIiIiZmZmIiIiZmZmZmZmZmZmZmZmZmZmIiIiIiIh3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERERERERERERERERERVVVVVVVVVVVVERERERERERERERERERERERERVVVVVVVVmZmZ3d3eIiIiIiIiIiIh3d3dmZmZEREREREREREQzMzNEREREREQzMzNEREREREQzMzMzMzMzMzMiIiIzMzMiIiIA//8AADMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzM0RERFVVVVVVVURERERERDMzMzMzM0RERERERERERDMzMyIiIjMzMzMzMyIiIjMzMyIiIjMzMzMzM0RERDMzMyIiIjMzMyIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERERERERERFVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVWZmZlVVVURERERERERERDMzM1VVVVVVVVVVVVVVVWZmZlVVVVVVVWZmZmZmZmZmZmZmZmZmZkRERDMzMzMzM0RERERERERERERERDMzM0RERERERDMzMzMzMzMzMzMzMzMzM0RERDMzMyIiIjMzMyIiIjMzMzMzM0RERERERERERERERDMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzM0RERGZmZlVVVTMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMyIiIjMzM0RERDMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIhERERERESIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzM0RERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVWZmZmZmZmZmZmZmZlVVVURERERERERERERERFVVVWZmZmZmZkRERERERERERERERERERERERERERFVVVVVVVURERFVVVURERERERERERDMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERDMzMzMzMyIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzM0RERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERERERERERERERDMzM0RERDMzM0RERERERDMzM0RERERERERERDMzM0RERERERFVVVURERERERDMzMzMzMzMzMyIiIjMzMzMzM0RERCIiIjMzMzMzMyIiIjMzMyIiIjMzMzMzMyIiIjMzMyIiIjMzM0RERERERFVVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERERERERERERERERERERERDMzMzMzM0RERERERERERFVVVURERERERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVURERERERDMzMzMzMzMzMzMzM0RERFVVVVVVVVVVVURERERERERERERERDMzM0RERERERERERFVVVVVVVWZmZmZmZnd3d2ZmZmZmZlVVVURERERERGZmZmZmZlVVVURERERERFVVVURERDMzM0RERERERERERERERERERFVVVURERERERERERFVVVVVVVVVVVVVVVURERERERERERERERDMzMzMzMzMzMzMzM0RERDMzMzMzM0RERDMzMzMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzM1VVVURERDMzMzMzMzMzMyIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzM0RERERERERERDMzMzMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIjMzMyIiIiIiIhERESIiIhERESIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzM0RERDMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMxERESIiIiIiIiIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIhERERERERERESIiIiIiIhERERERESIiIhERESIiIhERESIiIhERESIiIiIiIiIiIjMzMyIiIiIiIkRERDMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVVVVVWZmZnd3d3d3d3d3d4iIiJmZmaqqqszMzO7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7////////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7////u7u7u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7MzMzMzMzMzMzd3d3d3d3u7u7u7u7u7u7u7u7u7u7////u7u7u7u7d3d3d3d3MzMy7u7uqqqqZmZmZmZmIiIiZmZmZmZmIiIh3d3eIiIhmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3eIiIiIiIiIiIiIiIh3d3eIiIiIiIh3d3d3d3dmZmZ3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVEREQzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzNERERERERVVVVVVVVmZmZ3d3d3d3eIiIh3d3eIiIiIiIiIiIiZmZmZmZmIiIh3d3dmZmZmZmZmZmZVVVVERERERERERERERERERERERERERERERERERERERERVVVVVVVVVVVVmZmZmZmZVVVVVVVVEREREREREREREREQzMzNEREREREREREREREREREQzMzNEREQzMzNERERVVVVVVVWIiIh3d3eIiIh3d3dVVVUzMzNERERVVVVEREREREQzMzMzMzMzMzMzMzNEREQzMzNVVVUzMzMzMzMiIiIzMzMiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzNEREQzMzNERERVVVVEREQzMzMzMzNEREREREQzMzMzMzMzMzMiIiIzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzNEREQzMzNERERERERVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVEREREREQzMzNERERERERERERVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVEREREREQzMzMzMzNEREREREQzMzMzMzNEREREREQzMzMiIiIzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMiIiIzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIiIiIiIiIREREiIiIzMzMzMzMzMzMzMzMiIiIzMzMzMzNERERVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNEREQzMzMzMzMzMzMzMzNEREREREQzMzMiIiIiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIzMzNEREQzMzMiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzNVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERERERERERVVVVVVVVEREREREREREQzMzMzMzMiIiJERERmZmZVVVVVVVVERERVVVVVVVVERERERERERERVVVVVVVVVVVVEREREREREREREREQzMzMzMzMzMzMiIiIzMzNEREREREREREREREREREQiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIREREiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREREREQzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzNEREREREREREREREQzMzNEREREREREREQzMzMzMzMzMzNEREREREREREREREQzMzNERERVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMiIiIzMzMiIiIiIiIiIiIzMzMzMzMzMzMzMzNERERERERERERVVVVmZmZmZmZVVVVERERVVVVVVVVVVVVERERVVVUzMzNEREREREREREREREREREQzMzMzMzMzMzMzMzMzMzNERERVVVVERERERERVVVVmZmZERERERERVVVVERERVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVEREREREREREQzMzMzMzNERERERERERERERERVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERERERERERERERVVVVVVVVVVVVERERVVVV3d3d3d3dmZmZVVVVVVVVERERERERVVVVERERVVVVERERVVVVVVVVVVVVERERERERVVVVmZmZmZmZEREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMiIiIzMzNEREQzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzMiIiIzMzMiIiIzMzNEREREREREREREREREREREREREREQzMzNEREREREQzMzMzMzNEREREREQzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIzMzMiIiIiIiIREREREREiIiIREREiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIREREiIiIREREiIiIREREiIiIREREiIiIREREiIiIiIiIREREiIiIREREiIiIREREiIiIREREiIiIREREREREiIiIREREREREiIiIiIiIiIiIiIiIiIiIzMzMiIiJEREQzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzNERERERERVVVVVVVVmZmZmZmZ3d3eIiIiIiIiZmZnMzMzd3d3///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3dzMzM3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzM3d3d3d3d3d3dzMzM3d3dzMzM3d3d3d3d3d3d3d3d3d3dzMzM3d3d3d3d3d3d3d3dzMzMzMzM3d3d3d3d3d3d3d3d7u7u3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u////7u7u////////7u7u////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3d3d3d3d3d7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3dzMzMu7u7mZmZiIiId3d3d3d3d3d3ZmZmZmZmVVVVZmZmVVVVZmZmZmZmVVVVZmZmZmZmVVVVZmZmZmZmZmZmVVVVVVVVZmZmZmZmd3d3ZmZmZmZmZmZmd3d3iIiId3d3ZmZmZmZmd3d3ZmZmd3d3VVVVVVVVREREVVVVREREREREREREREREREREREREMzMzMzMzMzMzREREREREMzMzMzMzMzMzMzMzREREMzMzREREREREREREVVVVZmZmd3d3d3d3iIiIiIiId3d3d3d3d3d3iIiIiIiIiIiId3d3d3d3ZmZmd3d3ZmZmVVVVREREREREREREVVVVREREREREREREVVVVMzMzREREREREREREREREREREVVVVREREREREREREREREREREMzMzMzMzMzMzREREREREREREREREMzMzMzMzREREREREVVVVZmZmVVVVZmZmZmZmREREREREMzMzREREMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzREREREREREREREREREREREREMzMzMzMzMzMzREREMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzREREREREREREREREREREVVVVVVVVZmZmVVVVREREREREREREREREREREREREREREREREVVVVREREREREVVVVVVVVREREVVVVZmZmVVVVVVVVVVVVVVVVREREREREREREVVVVVVVVMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiMzMzIiIiMzMzMzMzREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzMzMzMzMzREREREREMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzIiIiMzMzREREREREVVVVVVVVREREREREMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREMzMzMzMzMzMzREREMzMzREREMzMzMzMzMzMzREREVVVVVVVVREREVVVVREREREREVVVVREREREREREREREREREREREREREREREREREREREREREREMzMzMzMzMzMzREREVVVVMzMzMzMzMzMzIiIiIiIiERERERERERERIiIiIiIiERERIiIiERERIiIiIiIiIiIiMzMzMzMzIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREMzMzREREREREREREMzMzIiIiMzMzREREMzMzMzMzMzMzREREMzMzREREMzMzREREREREREREMzMzREREREREREREREREREREREREREREVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiMzMzMzMzMzMzREREREREREREREREVVVVd3d3ZmZmVVVVVVVVVVVVVVVVREREREREREREREREMzMzREREREREREREREREMzMzMzMzMzMzREREREREREREREREREREVVVVVVVVVVVVVVVVREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVREREVVVVREREMzMzMzMzMzMzREREVVVVVVVVREREVVVVVVVVREREREREREREREREREREREREMzMzMzMzREREMzMzMzMzREREREREREREMzMzREREREREVVVVREREREREREREVVVVd3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREZmZmZmZmVVVVMzMzREREMzMzREREMzMzMzMzREREREREREREREREMzMzMzMzMzMzREREREREMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzREREVVVVREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzMzMzIiIiIiIiMzMzIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzREREMzMzIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiERERIiIiIiIiERERIiIiERERIiIiIiIiIiIiERERIiIiIiIiIiIiERERERERIiIiIiIiERERERERERERIiIiERERIiIiIiIiERERERERIiIiIiIiMzMzIiIiIiIiREREREREMzMzIiIiIiIiIiIiMzMzIiIiIiIiMzMzMzMzMzMzREREREREREREVVVVVVVVZmZmZmZmd3d3iIiIiIiImZmZzMzM7u7u////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////+7u7v///////+7u7v///+7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3czMzMzMzMzMzLu7u7u7u7u7u8zMzMzMzMzMzMzMzN3d3czMzMzMzMzMzMzMzMzMzMzMzLu7u8zMzMzMzLu7u7u7u8zMzMzMzMzMzLu7u7u7u7u7u7u7u8zMzMzMzMzMzMzMzMzMzMzMzMzMzN3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3d3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////+7u7v///////////////////////////+7u7v///////////////////+7u7v///////////////////////////////////////+7u7u7u7u7u7t3d3e7u7u7u7v///+7u7v///+7u7u7u7v///+7u7u7u7t3d3czMzKqqqoiIiHd3d2ZmZmZmZlVVVVVVVURERERERERERERERERERERERFVVVURERFVVVURERFVVVVVVVURERFVVVVVVVURERGZmZlVVVVVVVWZmZmZmZnd3d3d3d3d3d3d3d4iIiHd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d1VVVVVVVURERERERERERERERDMzM0RERDMzM0RERERERERERDMzM0RERERERDMzM0RERERERFVVVXd3d3d3d4iIiHd3d4iIiHd3d3d3d2ZmZnd3d2ZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZlVVVURERFVVVVVVVVVVVWZmZkRERERERERERERERERERDMzM0RERERERERERERERFVVVWZmZlVVVVVVVURERERERDMzM0RERERERERERDMzMzMzMzMzMzMzM0RERFVVVURERERERERERERERDMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzM0RERERERDMzM0RERERERDMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzM0RERERERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzM0RERDMzM0RERERERERERERERERERFVVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERERERERERFVVVURERERERFVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERFVVVURERERERDMzMzMzM0RERERERERERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzM0RERERERERERCIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzM0RERERERERERDMzMzMzM0RERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERDMzM0RERERERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERFVVVVVVVVVVVURERDMzMzMzMzMzM0RERFVVVWZmZmZmZkRERERERDMzMzMzMzMzM0RERERERERERERERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVURERERERFVVVURERERERFVVVURERERERERERERERERERDMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERFVVVTMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIjMzM0RERDMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERERERERERDMzMzMzMzMzM0RERERERERERFVVVTMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM0RERDMzMzMzM0RERERERERERERERFVVVVVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzM0RERERERERERERERERERERERGZmZmZmZlVVVVVVVWZmZlVVVURERDMzM0RERERERERERDMzM0RERERERDMzM0RERERERERERERERERERDMzM0RERDMzM1VVVVVVVVVVVVVVVURERERERERERERERERERFVVVVVVVVVVVVVVVURERFVVVURERDMzMzMzMzMzM0RERFVVVURERERERFVVVVVVVURERERERDMzM0RERDMzMzMzM0RERDMzMzMzMzMzM0RERERERERERCIiIjMzMzMzMzMzMzMzM0RERERERDMzM1VVVWZmZnd3d2ZmZlVVVWZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d2ZmZlVVVURERERERFVVVWZmZlVVVURERERERERERERERERERERERDMzM0RERERERERERERERERERERERDMzM0RERFVVVTMzMyIiIjMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERERERDMzMzMzM0RERERERERERERERERERERERERERERERDMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzMyIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIjMzMyIiIiIiIjMzMyIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIjMzM0RERERERDMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzMyIiIjMzMyIiIhERESIiIhERERERESIiIhERESIiIhERERERESIiIiIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzM0RERDMzMyIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzM0RERERERERERFVVVWZmZnd3d3d3d4iIiJmZmaqqqszMzN3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////u7u7////////////////////////////////////////u7u7u7u7u7u7d3d3u7u7u7u7u7u7d3d3u7u7d3d3d3d3MzMzMzMy7u7u7u7u7u7vMzMzMzMzd3d3MzMzd3d3d3d3d3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMy7u7vMzMy7u7vMzMy7u7vMzMy7u7u7u7u7u7u7u7u7u7u7u7u7u7uqqqq7u7u7u7vMzMy7u7vMzMzMzMzMzMzMzMzd3d3d3d3MzMzd3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7////u7u7////////////u7u7////////u7u7////////u7u7////////u7u7////////////////////////////////u7u7////////u7u7////////u7u7////////////u7u7////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7d3d3u7u7u7u7u7u7u7u7u7u7////////u7u7u7u7u7u7u7u7d3d27u7uZmZmIiIh3d3dmZmZmZmZERERVVVVVVVVVVVVERERERERVVVVERERVVVVERERERERERERERERERERERERVVVVERERVVVVVVVVVVVVVVVVmZmZmZmaIiIiIiIiIiIiZmZmIiIh3d3eIiIiIiIiIiIiZmZmIiIiZmZmqqqqIiIhmZmZ3d3d3d3dVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVERERERERVVVVmZmZ3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3d3d3dmZmZmZmZ3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVEREREREREREQzMzNERERVVVVVVVVmZmZmZmZmZmZmZmZ3d3d3d3dmZmZVVVVVVVUzMzMzMzMiIiIzMzMzMzMzMzMzMzNEREQzMzNEREQzMzNEREQzMzMzMzMiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIzMzMzMzMzMzNERERERERVVVVEREREREQzMzMzMzMzMzMzMzNEREQiIiIiIiIzMzMiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIzMzMiIiIiIiIzMzMzMzMzMzNEREQzMzMzMzNERERERERERERVVVVERERVVVVERERERERVVVVVVVVERERVVVVEREQzMzNVVVVERERERERERERERERVVVVERERVVVVmZmZVVVVVVVVEREREREQzMzNERERERERVVVVEREREREREREREREQzMzNEREQzMzMzMzMzMzMiIiIzMzNEREREREREREQzMzMzMzMzMzMiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzMiIiIiIiIzMzMzMzNEREREREREREREREREREREREQzMzNVVVVEREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzNEREQzMzNEREQzMzNEREREREQzMzNEREQzMzNEREQzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMiIiIzMzNERERERERVVVVERERERERERERERERVVVVEREREREREREQzMzNEREQzMzMiIiIzMzNVVVVmZmZEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERERERERERERERVVVVVVVVEREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzNEREREREQzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiJERERVVVVEREQiIiIzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNVVVVEREREREQzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzNEREQzMzMzMzMzMzNERERERERERERERERERERVVVVmZmZVVVVEREQzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzNERERERERERERERERERERERERmZmZ3d3dVVVVmZmZVVVVVVVVVVVVEREREREREREQzMzMzMzNEREQzMzNEREQzMzNERERERERERERVVVVERERERERVVVVVVVVERERERERVVVVERERERERERERERERERERVVVVERERVVVVERERERERERERERERERERERERERERERERERERERERVVVVmZmZVVVVEREREREREREQzMzMzMzNEREREREQzMzNEREQzMzNEREQzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNERERmZmZmZmZERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3eIiIh3d3dmZmZVVVVVVVVmZmZmZmZVVVVEREREREQzMzNEREQzMzNEREQzMzNEREREREREREREREREREREREQzMzNVVVVEREQzMzMzMzNEREQzMzMiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMiIiIzMzMzMzNEREREREQzMzMzMzNEREREREREREREREQzMzNEREQzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVEREQiIiIzMzMiIiIzMzMiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIREREiIiIiIiIiIiIREREREREiIiIiIiIiIiIzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIREREiIiIiIiIREREiIiIREREiIiIiIiIREREREREiIiIREREiIiIiIiIzMzMzMzMiIiIiIiIREREiIiIREREREREREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiJEREQzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzMzMzNERERERERERERVVVVVVVVmZmZ3d3d3d3eZmZmqqqq7u7vd3d3u7u7u7u7////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM3d3d3d3d3d3dzMzMzMzMzMzM3d3dzMzM3d3dzMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7qqqqu7u7u7u7u7u7qqqqu7u7qqqqu7u7u7u7zMzMzMzMzMzM3d3d3d3d3d3d3d3dzMzMzMzM3d3dzMzMzMzMzMzMzMzM3d3d3d3d7u7u7u7u7u7u7u7u////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////7u7u////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u////////7u7u7u7u////7u7u7u7u7u7uzMzMzMzMqqqqiIiId3d3d3d3VVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiImZmZmZmZmZmZqqqqqqqqqqqqu7u7qqqqmZmZd3d3d3d3d3d3ZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmVVVVZmZmVVVVVVVVd3d3ZmZmd3d3ZmZmd3d3ZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVREREREREVVVVREREREREREREREREREREREREREREREREVVVVREREREREVVVVREREREREREREVVVVZmZmZmZmd3d3iIiImZmZiIiIVVVVREREMzMzMzMzMzMzMzMzREREMzMzMzMzREREREREREREMzMzMzMzIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzMzMzREREMzMzREREREREREREREREMzMzMzMzIiIiMzMzREREMzMzIiIiMzMzIiIiIiIiIiIiMzMzIiIiIiIiMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzMzMzREREREREREREREREREREVVVVREREVVVVVVVVREREREREREREREREREREREREVVVVREREREREREREREREVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREMzMzREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREMzMzMzMzMzMzIiIiMzMzMzMzIiIiMzMzMzMzMzMzREREMzMzMzMzREREREREMzMzMzMzIiIiMzMzMzMzIiIiMzMzMzMzIiIiMzMzREREREREREREREREREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREMzMzREREMzMzMzMzMzMzREREZmZmREREREREMzMzMzMzREREMzMzREREREREREREREREMzMzREREMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzIiIiIiIiREREREREREREREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiREREREREREREREREREREMzMzREREMzMzREREREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzREREREREMzMzREREMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzREREREREMzMzIiIiIiIiIiIiMzMzREREMzMzMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREREREMzMzREREMzMzMzMzMzMzREREREREMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREMzMzREREREREREREREREREREVVVVVVVVVVVVMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzREREREREVVVVVVVVREREZmZmd3d3ZmZmVVVVZmZmZmZmVVVVVVVVMzMzMzMzMzMzMzMzREREREREMzMzREREREREMzMzREREREREREREREREREREREREVVVVZmZmREREREREREREREREREREREREREREREREREREREREREREREREREREREREMzMzREREREREREREMzMzREREVVVVVVVVREREREREMzMzREREMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREMzMzREREREREREREREREREREREREREREMzMzREREREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3ZmZmREREVVVVZmZmZmZmVVVVREREMzMzMzMzMzMzREREREREREREREREREREZmZmVVVVREREMzMzREREREREREREMzMzREREMzMzIiIiIiIiIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREREREMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREREREMzMzREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzIiIiIiIiERERERERERERIiIiIiIiERERIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzIiIiERERERERIiIiIiIiIiIiIiIiERERERERIiIiIiIiIiIiIiIiIiIiERERIiIiMzMzIiIiMzMzIiIiIiIiERERIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzREREREREREREREREVVVVZmZmd3d3iIiImZmZqqqqzMzM3d3d7u7u7u7u////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////+7u7v///////////////////////////////////+7u7v///////+7u7u7u7u7u7t3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3czMzMzMzN3d3d3d3e7u7t3d3d3d3d3d3czMzN3d3d3d3czMzMzMzLu7u8zMzLu7u8zMzLu7u7u7u7u7u7u7u6qqqru7u7u7u7u7u7u7u8zMzMzMzN3d3czMzN3d3d3d3czMzMzMzMzMzN3d3czMzMzMzMzMzMzMzN3d3d3d3d3d3e7u7u7u7u7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////+7u7v///+7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3e7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7v///+7u7u7u7u7u7u7u7v///+7u7v///+7u7u7u7u7u7u7u7u7u7v///+7u7v///////+7u7v///+7u7u7u7t3d3czMzKqqqpmZmXd3d3d3d2ZmZmZmZlVVVWZmZlVVVWZmZmZmZnd3d3d3d2ZmZnd3d2ZmZmZmZlVVVVVVVURERFVVVVVVVXd3d4iIiIiIiHd3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d3d3d3d3d4iIiIiIiJmZmZmZmaqqqpmZmaqqqpmZmaqqqoiIiHd3d3d3d2ZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVWZmZmZmZmZmZlVVVVVVVWZmZnd3d3d3d4iIiHd3d4iIiHd3d2ZmZnd3d3d3d2ZmZmZmZnd3d1VVVVVVVURERFVVVURERERERERERERERFVVVURERERERDMzM0RERERERERERERERERERFVVVURERERERERERFVVVWZmZnd3d3d3d4iIiKqqqqqqqmZmZkRERERERDMzMzMzM0RERDMzMzMzMzMzMzMzM0RERERERDMzMyIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIjMzMzMzMyIiIiIiIjMzMzMzMzMzMyIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzM0RERERERDMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzM0RERDMzMyIiIjMzMzMzMzMzMzMzM0RERERERFVVVURERERERERERFVVVVVVVVVVVURERERERERERERERERERERERERERFVVVURERERERERERFVVVVVVVURERFVVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVURERERERDMzMzMzMzMzMzMzM0RERERERERERERERDMzMzMzMzMzM0RERFVVVURERERERDMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERERERDMzMzMzMzMzMzMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERERERERERFVVVURERERERFVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERDMzM0RERERERDMzMzMzMzMzM0RERGZmZlVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzM0RERFVVVURERERERDMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERERERERERDMzM0RERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIjMzM0RERERERDMzMzMzMzMzMyIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzM1VVVURERDMzMyIiIjMzMzMzM0RERERERERERDMzM0RERDMzMzMzMzMzM0RERDMzMzMzMzMzM0RERDMzM0RERDMzMzMzMzMzM0RERERERERERDMzMzMzMzMzM0RERDMzM0RERERERDMzMzMzMyIiIjMzMyIiIjMzM0RERERERERERERERERERERERERERFVVVVVVVWZmZkRERDMzMzMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERFVVVURERERERFVVVVVVVWZmZnd3d1VVVWZmZmZmZmZmZkRERERERDMzMzMzMzMzMzMzM0RERERERERERERERERERERERERERERERERERERERFVVVVVVVVVVVURERERERERERERERFVVVURERFVVVURERERERERERERERERERERERDMzM0RERERERERERERERERERERERFVVVVVVVVVVVURERERERDMzM0RERERERDMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERERERERERERERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVURERGZmZnd3d2ZmZlVVVURERERERERERDMzM0RERERERERERERERFVVVVVVVURERDMzMzMzM0RERERERFVVVTMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERDMzMzMzM0RERDMzMzMzMzMzM0RERERERERERERERDMzM0RERFVVVVVVVURERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERDMzMyIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIhERESIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzM0RERDMzMzMzMzMzMyIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIhERESIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzM0RERDMzMzMzMzMzM0RERDMzMyIiIjMzMyIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzM0RERERERERERFVVVWZmZmZmZoiIiJmZmbu7u8zMzN3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3d3d3d3d3d3d3d3d3u7u7d3d3d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7uqqqq7u7uqqqrMzMy7u7u7u7vMzMzd3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzd3d3d3d3d3d3MzMzd3d3u7u7d3d3u7u7////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////d3d3d3d3MzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7vMzMzMzMzMzMzd3d3MzMzd3d3d3d3d3d3MzMzd3d3MzMzMzMy7u7u7u7vMzMy7u7vd3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzd3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7////u7u7u7u7u7u7u7u7u7u7d3d3d3d3MzMyqqqqqqqqIiIiIiIh3d3dmZmZmZmZVVVVVVVVVVVVmZmZ3d3d3d3d3d3dmZmZmZmZmZmZVVVVVVVVVVVVmZmZ3d3eIiIiZmZmZmZmIiIiIiIiIiIiIiIiIiIh3d3dmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3eIiIiIiIh3d3eIiIiZmZmIiIh3d3d3d3d3d3eIiIiIiIh3d3dmZmZmZmZVVVVmZmZmZmZ3d3d3d3d3d3dmZmZmZmZmZmZ3d3d3d3eIiIiIiIiIiIiIiIh3d3d3d3dmZmZ3d3dmZmZmZmZERERVVVVEREREREQzMzMzMzMzMzNEREQzMzMzMzNEREQzMzNEREREREREREREREQzMzNEREREREREREQzMzNERERmZmZ3d3dmZmaIiIiZmZl3d3dVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzNEREQiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzMiIiIzMzMiIiJEREQzMzMiIiIiIiIzMzNEREQzMzNERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVERERERERERERERERVVVVEREREREQzMzNVVVVERERERERERERERERERERVVVVVVVVERERERERERERERERVVVVVVVVEREREREQzMzNEREREREREREQzMzNERERVVVVEREQzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMiIiIiIiIiIiIzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREREREREREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERERERVVVVVVVVVVVVVVVVEREQzMzMzMzNERERVVVVmZmZVVVUzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIiIiIzMzMiIiIzMzNEREREREREREREREREREQzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzNEREQzMzMzMzNEREREREREREQzMzNERERVVVVEREREREREREREREREREREREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIzMzMzMzNERERVVVUzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzNVVVVmZmZEREQzMzMzMzMzMzMiIiIzMzMzMzNEREREREQzMzNEREQzMzNEREQzMzNEREQzMzNEREREREQzMzNEREQzMzNERERERERVVVVVVVVEREQzMzMzMzNEREREREREREQzMzMzMzMiIiIzMzMzMzMzMzMzMzNERERERERERERERERERERVVVVERERERERmZmZVVVVEREQzMzMiIiIiIiIzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzNERERERERVVVVERERVVVVERERVVVVVVVVERERVVVVVVVVVVVV3d3dmZmZmZmZEREQzMzMzMzNEREQzMzNERERERERVVVVERERERERVVVVERERERERERERVVVVERERVVVVVVVVERERERERVVVVERERVVVVERERVVVVEREREREREREREREREREQzMzNEREQzMzNEREREREREREQzMzNERERVVVVERERVVVVVVVVVVVVEREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzNERERERERERERERERVVVVERERERERVVVVERERERERERERERERVVVVERERVVVVERERVVVVmZmZmZmZVVVVmZmZmZmZVVVVERERVVVVERERVVVVVVVVmZmZVVVVVVVUzMzMzMzMzMzNVVVVmZmZEREQzMzMzMzMiIiIzMzNEREREREREREREREQzMzMzMzMiIiIzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzNERERERERERERERERERERERERERERERERVVVVVVVVEREREREREREQzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNEREQzMzMiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIzMzNEREREREREREQzMzMiIiIiIiIzMzMzMzNEREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzNERERVVVVmZmZmZmZ3d3eZmZm7u7vMzMzMzMzu7u7u7u7u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////7u7u3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7u7u7zMzMzMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7zMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d7u7u3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzM3d3dzMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7zMzMzMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3dzMzMzMzMu7u7zMzMzMzMu7u7zMzMzMzM3d3d3d3d7u7u7u7u7u7u////7u7u////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3dzMzMzMzMzMzMu7u7zMzMzMzMu7u7u7u7zMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzM3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3d3d3dzMzMzMzMu7u7u7u7u7u7zMzMzMzMzMzM7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3dzMzMzMzMu7u7u7u7qqqqmZmZqqqqiIiId3d3d3d3ZmZmZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVZmZmiIiImZmZiIiIiIiIiIiIiIiIiIiId3d3ZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmd3d3d3d3iIiIiIiIiIiId3d3d3d3ZmZmd3d3d3d3ZmZmVVVVVVVVVVVVVVVVVVVVZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmVVVVVVVVREREREREREREREREMzMzMzMzIiIiMzMzREREREREIiIiMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzMzMzMzMzREREREREREREVVVVZmZmd3d3VVVVMzMzMzMzMzMzIiIiIiIiMzMzMzMzMzMzMzMzIiIiERERERERIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzIiIiIiIiMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzREREREREVVVVVVVVREREREREREREVVVVVVVVREREREREREREREREVVVVREREREREMzMzREREREREREREREREREREREREREREREREREREMzMzMzMzREREMzMzREREVVVVVVVVREREREREMzMzREREREREREREREREVVVVVVVVMzMzREREMzMzMzMzREREREREMzMzMzMzMzMzMzMzREREREREMzMzMzMzIiIiMzMzMzMzIiIiMzMzMzMzMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREREREREREREREREREREREMzMzREREREREREREMzMzREREMzMzMzMzREREMzMzMzMzREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVREREMzMzMzMzMzMzMzMzVVVVVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzREREREREREREMzMzMzMzMzMzMzMzREREVVVVVVVVREREREREREREMzMzREREREREMzMzREREREREREREREREMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzMzMzIiIiMzMzREREVVVVREREREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzVVVVVVVVREREMzMzMzMzIiIiMzMzREREMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREREREREREMzMzVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzREREMzMzMzMzMzMzREREREREREREREREREREVVVVVVVVZmZmZmZmREREMzMzIiIiMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzREREVVVVREREVVVVVVVVREREVVVVREREVVVVVVVVREREREREVVVVd3d3VVVVREREMzMzMzMzREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVREREREREREREREREVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREREREREREREREREREREREREREMzMzREREREREVVVVREREREREREREVVVVVVVVREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVVVVVREREREREREREMzMzREREREREREREVVVVVVVVREREVVVVREREREREREREMzMzREREREREVVVVMzMzVVVVVVVVVVVVd3d3d3d3ZmZmVVVVZmZmVVVVZmZmZmZmd3d3d3d3d3d3VVVVREREMzMzVVVViIiIZmZmREREMzMzREREMzMzREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREMzMzREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVREREREREREREREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzREREMzMzREREMzMzMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzMzMzIiIiMzMzIiIiERERIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiERERIiIiIiIiMzMzVVVVVVVVREREMzMzREREREREMzMzREREMzMzMzMzIiIiREREMzMzREREMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzREREREREVVVVVVVVd3d3mZmZqqqqu7u7zMzM3d3d7u7u7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////+7u7v///////////////////+7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u7u7u6qqqqqqqru7u7u7u7u7u7u7u8zMzN3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzN3d3czMzN3d3d3d3d3d3czMzN3d3czMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u8zMzLu7u93d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3czMzMzMzLu7u7u7u7u7u8zMzMzMzMzMzN3d3d3d3e7u7u7u7u7u7v///////////////////+7u7v///////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////+7u7u7u7u7u7u7u7u7u7t3d3d3d3czMzMzMzMzMzN3d3czMzN3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzN3d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzLu7u7u7u7u7u7u7u6qqqru7u7u7u6qqqpmZmZmZmYiIiIiIiIiIiHd3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZnd3d3d3d4iIiIiIiIiIiIiIiJmZmXd3d2ZmZmZmZlVVVWZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiIiIiHd3d3d3d4iIiHd3d2ZmZlVVVWZmZlVVVURERERERERERERERERERERERFVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVXd3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVURERERERERERDMzMzMzM0RERERERERERCIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERDMzM0RERDMzMzMzM0RERERERERERERERDMzMzMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzM0RERFVVVURERERERERERERERERERERERERERERERDMzMzMzM0RERFVVVURERERERDMzM0RERERERERERERERERERDMzM0RERERERERERERERDMzM0RERDMzM0RERERERFVVVURERERERDMzM0RERERERDMzMzMzM0RERFVVVVVVVTMzM0RERERERERERERERDMzM0RERDMzM0RERDMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzM0RERERERDMzM0RERDMzM0RERERERERERERERERERERERERERERERERERFVVVURERERERERERERERDMzM0RERFVVVURERERERERERDMzM0RERDMzM1VVVURERFVVVWZmZmZmZlVVVVVVVVVVVURERFVVVTMzMzMzMzMzMyIiIjMzM0RERERERERERDMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMzMzMyIiIjMzMyIiIiIiIiIiIjMzMzMzMyIiIjMzM0RERERERFVVVURERDMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERDMzMzMzMzMzM0RERERERFVVVWZmZlVVVURERDMzM0RERERERDMzMzMzM0RERFVVVURERERERDMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzM0RERERERFVVVVVVVWZmZlVVVTMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIjMzMyIiIjMzMzMzMyIiIjMzMyIiIiIiIjMzM1VVVURERDMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERERERDMzMzMzMzMzMzMzM0RERERERDMzM0RERERERERERERERDMzMzMzM0RERERERERERDMzM0RERDMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERERERERERERERERERFVVVXd3d2ZmZlVVVVVVVTMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERERERFVVVVVVVURERERERFVVVURERFVVVURERFVVVURERERERERERERERERERDMzMzMzM0RERERERERERERERERERERERFVVVVVVVVVVVVVVVURERFVVVURERERERERERFVVVVVVVVVVVVVVVVVVVURERERERDMzM0RERDMzM0RERDMzM0RERERERERERERERERERERERERERERERERERERERFVVVVVVVVVVVVVVVURERERERDMzM0RERDMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM0RERDMzM0RERGZmZmZmZlVVVURERDMzM0RERERERDMzM0RERFVVVURERERERERERERERERERERERERERDMzM0RERERERERERERERERERFVVVWZmZnd3d2ZmZmZmZlVVVVVVVVVVVVVVVWZmZnd3d4iIiHd3d2ZmZkRERFVVVXd3d2ZmZlVVVVVVVURERERERDMzM0RERERERERERDMzM0RERERERERERDMzM0RERERERDMzM0RERERERDMzMzMzMzMzM1VVVVVVVURERFVVVURERFVVVWZmZlVVVVVVVVVVVVVVVURERDMzM0RERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERDMzMzMzMyIiIiIiIiIiIjMzM0RERDMzMzMzMzMzMyIiIiIiIjMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzM0RERDMzMzMzMzMzMyIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIhERESIiIiIiIhERESIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzM0RERFVVVURERERERERERDMzMzMzMzMzMyIiIjMzMzMzM0RERDMzM0RERDMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIhERESIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIkRERERERERERFVVVXd3d4iIiJmZmaqqqru7u8zMzN3d3e7u7u7u7v///////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////u7u7////////////////////u7u7////////u7u7u7u7u7u7u7u7u7u7d3d3d3d3MzMzMzMzMzMzMzMy7u7u7u7uqqqq7u7uqqqq7u7u7u7u7u7u7u7u7u7vMzMzMzMzd3d3MzMy7u7vMzMy7u7vMzMzMzMzMzMzMzMzd3d3MzMzd3d3MzMzMzMzd3d3MzMzd3d3d3d3d3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3d3d3d3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMzMzMy7u7uqqqqqqqqqqqq7u7u7u7u7u7u7u7vMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMy7u7vMzMy7u7u7u7vMzMzd3d3d3d3u7u7u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3d3d3d3d3u7u7d3d3u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzd3d3d3d3MzMzd3d3MzMzMzMzMzMzMzMzMzMzd3d3d3d3d3d3u7u7d3d3d3d3d3d3d3d3d3d3MzMzd3d3MzMy7u7u7u7u7u7uZmZmqqqqqqqqqqqqqqqqZmZmZmZmZmZmZmZmIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3dmZmZmZmZmZmaIiIh3d3eIiIiZmZmZmZmZmZmZmZmIiIh3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3eIiIiIiIiIiIiIiIh3d3dVVVVEREREREREREREREREREREREQzMzMzMzMzMzNERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZEREREREQzMzNERERVVVVVVVVVVVVmZmZ3d3d3d3dmZmZ3d3dVVVVEREQzMzMzMzNEREQzMzNEREQzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMREREiIiIREREREREiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzNEREREREQiIiIzMzMzMzNEREQzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMiIiIzMzMzMzNEREQzMzMzMzNEREREREREREREREREREREREREREREREQzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzNERERERERERERERERERERERERVVVVEREREREQzMzMzMzMzMzMzMzNERERmZmZVVVVERERVVVVEREREREQzMzMiIiJERERVVVVVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREREREREREREREQzMzNERERERERERERERERVVVVmZmZmZmZmZmZVVVUzMzNERERERERmZmZVVVVmZmZVVVVERERERERERERERERERERVVVVmZmZVVVVVVVVVVVVEREREREREREREREQzMzMzMzMzMzMzMzNVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzNEREQzMzNEREREREREREREREQzMzNVVVVmZmZVVVVEREREREQzMzNEREQzMzNEREREREREREREREREREQzMzMzMzMiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzNVVVVVVVVVVVVVVVVmZmZVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzMiIiIiIiJERERERERVVVVEREQzMzMzMzNEREREREQzMzMzMzMzMzNEREREREQzMzNEREQzMzMzMzNERERERERERERVVVVVVVVEREQzMzMzMzNEREREREREREREREQzMzMzMzMzMzMzMzNEREQzMzNEREREREQzMzMzMzNERERERERERERVVVVmZmZ3d3d3d3dmZmZERERVVVVEREREREQzMzNEREQzMzMzMzMzMzMiIiIzMzMzMzNERERERERERERERERERERVVVVERERERERVVVVERERERERVVVVEREQiIiIzMzNERERERERERERERERERERERERVVVVERERVVVVVVVVVVVVmZmZVVVVVVVVERERVVVVVVVVVVVVERERVVVVVVVVERERVVVVVVVVVVVVEREREREREREREREQzMzNERERERERERERVVVVVVVVVVVVVVVVERERERERERERERERVVVVVVVVVVVVVVVVVVVVEREREREQzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzNEREQzMzNEREQzMzNERERmZmZmZmZERERVVVVERERERERVVVVEREREREREREREREREREREREREREQzMzNEREREREREREREREREREREREQzMzNVVVVmZmZmZmZVVVVVVVVERERVVVVVVVVVVVVmZmZmZmZmZmZ3d3dmZmZVVVVVVVVmZmZ3d3dmZmZVVVVEREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREQzMzMzMzMzMzNVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVEREREREREREREREREREREREREREREREQzMzMiIiIzMzMzMzNEREREREQzMzNEREQzMzMzMzMzMzMzMzMiIiIiIiIzMzMzMzMzMzMiIiIREREiIiIiIiIzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIiIiIzMzMzMzNEREQzMzNEREREREREREREREQzMzMzMzMzMzMiIiIzMzMzMzNEREREREQzMzMzMzMzMzMzMzMiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIREREiIiIREREiIiIiIiIREREiIiIiIiIiIiIiIiIzMzNERERVVVVmZmZ3d3eIiIiqqqqqqqq7u7vMzMzd3d3d3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7u7u7u7u7zMzMzMzMu7u7zMzMzMzM3d3dzMzMzMzM3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzM3d3dzMzMzMzM3d3d3d3d3d3d3d3dzMzMzMzMzMzMu7u7u7u7qqqqqqqqqqqqqqqqmZmZmZmZu7u7u7u7zMzMzMzMzMzM3d3d3d3d7u7u3d3d7u7u7u7u7u7u3d3dzMzMzMzMu7u7qqqqu7u7qqqqu7u7zMzM3d3d3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u3d3d7u7u3d3d3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3dzMzMu7u7u7u7qqqqqqqqqqqqmZmZqqqqmZmZmZmZmZmZiIiId3d3d3d3d3d3iIiId3d3ZmZmd3d3iIiId3d3d3d3iIiId3d3d3d3iIiIiIiIiIiImZmZqqqqqqqqmZmZqqqqmZmZiIiIiIiId3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3iIiIZmZmREREREREMzMzREREREREMzMzREREREREREREMzMzREREVVVVZmZmVVVVREREREREREREREREVVVVZmZmZmZmVVVVVVVVREREVVVVZmZmZmZmVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3qqqqqqqqqqqqiIiImZmZiIiIVVVVMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiERERIiIiMzMzIiIiIiIiERERIiIiIiIiERERIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREREREMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREREREREREREREREREMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVREREMzMzMzMzREREVVVVVVVVREREREREREREREREMzMzMzMzREREMzMzMzMzREREVVVVVVVVVVVVVVVVREREMzMzMzMzMzMzIiIiMzMzMzMzREREMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzREREREREMzMzREREREREREREREREREREREREREREREREMzMzVVVVVVVVVVVVZmZmZmZmd3d3iIiId3d3d3d3d3d3REREREREREREVVVVZmZmZmZmVVVVMzMzREREREREREREREREREREREREREREVVVVVVVVREREREREREREMzMzMzMzMzMzMzMzREREREREVVVVREREMzMzMzMzIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzVVVVVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREREREREREREREREREREREREREREREMzMzVVVVZmZmREREMzMzMzMzREREREREREREREREREREMzMzMzMzMzMzIiIiMzMzIiIiIiIiMzMzMzMzMzMzREREREREREREREREVVVVREREZmZmd3d3ZmZmREREMzMzREREMzMzMzMzMzMzMzMzREREMzMzIiIiMzMzIiIiMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzREREVVVVVVVVREREREREREREMzMzMzMzMzMzMzMzREREMzMzREREMzMzREREREREREREREREREREVVVVZmZmREREMzMzREREREREREREREREREREREREMzMzMzMzMzMzREREREREREREREREREREMzMzMzMzREREREREZmZmd3d3d3d3d3d3VVVVVVVVREREVVVVREREMzMzREREREREMzMzMzMzMzMzMzMzREREREREREREREREREREVVVVREREREREREREREREREREREREREREREREMzMzIiIiMzMzREREVVVVVVVVREREVVVVREREVVVVVVVVVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVREREREREVVVVVVVVREREMzMzMzMzREREREREVVVVVVVVREREREREVVVVREREREREVVVVREREREREREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREZmZmVVVVVVVVVVVVREREREREVVVVVVVVREREREREREREREREREREREREREREVVVVREREVVVVREREREREREREREREVVVVREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmd3d3ZmZmZmZmd3d3VVVVVVVVVVVVVVVVREREREREVVVVVVVVREREREREREREREREREREMzMzMzMzVVVVVVVVREREVVVVREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzVVVVVVVVMzMzREREREREMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiERERIiIiMzMzREREREREMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzREREMzMzREREMzMzIiIiMzMzIiIiMzMzIiIiIiIiMzMzIiIiIiIiIiIiMzMzIiIiMzMzMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiMzMzREREREREREREREREREREIiIiMzMzMzMzMzMzMzMzREREVVVVVVVVMzMzIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiERERIiIiERERIiIiIiIiIiIiMzMzMzMzREREZmZmd3d3mZmZmZmZqqqqqqqqu7u7zMzM3d3d3d3d3d3d////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////+7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3e7u7u7u7u7u7u7u7t3d3e7u7t3d3e7u7t3d3d3d3czMzN3d3czMzN3d3czMzMzMzMzMzLu7u6qqqru7u6qqqqqqqqqqqqqqqru7u7u7u7u7u8zMzLu7u8zMzMzMzMzMzMzMzN3d3czMzN3d3d3d3czMzMzMzN3d3czMzMzMzN3d3czMzN3d3czMzMzMzMzMzMzMzMzMzN3d3d3d3d3d3czMzMzMzMzMzMzMzLu7u6qqqqqqqqqqqqqqqru7u7u7u7u7u7u7u7u7u8zMzMzMzMzMzN3d3d3d3d3d3e7u7u7u7t3d3d3d3d3d3bu7u6qqqqqqqpmZmaqqqqqqqru7u8zMzMzMzN3d3e7u7u7u7u7u7u7u7v///////////////////+7u7v///////////////////////////////////////////////////+7u7v///////+7u7v///////////////////////+7u7v///////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7u7u7t3d3d3d3czMzMzMzMzMzMzMzN3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3czMzN3d3czMzMzMzMzMzMzMzLu7u7u7u7u7u6qqqqqqqqqqqpmZmYiIiIiIiJmZmYiIiIiIiHd3d5mZmYiIiHd3d4iIiIiIiHd3d4iIiIiIiJmZmZmZmZmZmZmZmaqqqpmZmZmZmaqqqqqqqpmZmZmZmYiIiIiIiIiIiJmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiHd3d1VVVURERERERDMzMzMzMzMzM0RERDMzM0RERERERERERERERERERERERERERERERERERERERERERERERERERFVVVVVVVURERFVVVURERGZmZmZmZkRERERERGZmZmZmZlVVVURERFVVVVVVVWZmZnd3d1VVVWZmZmZmZnd3d5mZmaqqqqqqqqqqqnd3d1VVVTMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMyIiIhERERERESIiIiIiIiIiIiIiIjMzMyIiIhERERERERERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzM0RERCIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIkRERDMzM0RERDMzMzMzMzMzMzMzMzMzM0RERDMzMyIiIjMzMzMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzM1VVVVVVVURERERERERERERERERERERERDMzMzMzM0RERERERDMzMzMzM0RERERERFVVVURERERERDMzM0RERFVVVVVVVVVVVURERERERERERDMzMzMzMzMzM0RERERERDMzM0RERERERFVVVURERERERERERDMzMyIiIiIiIhERETMzMzMzM0RERDMzMzMzMzMzMzMzM0RERFVVVURERERERERERDMzM0RERDMzMzMzM0RERERERDMzM0RERERERFVVVURERERERERERDMzMzMzM0RERERERFVVVWZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZlVVVVVVVURERERERERERGZmZlVVVURERERERFVVVURERERERERERERERFVVVURERFVVVVVVVVVVVURERERERDMzMzMzMzMzM0RERERERERERFVVVTMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERDMzM0RERDMzMzMzM0RERFVVVURERERERERERERERERERERERERERERERERERERERERERERERERERERERGZmZlVVVURERERERDMzM0RERERERERERDMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzM0RERERERERERERERDMzMzMzM0RERFVVVVVVVURERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzM0RERDMzMyIiIjMzM0RERERERERERGZmZlVVVURERERERDMzMzMzM0RERDMzM0RERERERERERERERERERERERERERERERERERERERERERFVVVURERERERERERERERERERERERERERDMzMzMzMzMzM1VVVURERERERERERERERERERDMzM0RERFVVVWZmZmZmZnd3d2ZmZmZmZlVVVVVVVURERERERERERDMzMzMzM0RERERERERERDMzM0RERERERDMzM0RERDMzM0RERERERERERDMzMzMzM0RERERERERERERERERERDMzMzMzM0RERERERFVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVURERERERERERERERERERERERDMzM0RERERERERERFVVVVVVVVVVVURERERERERERFVVVVVVVURERERERERERERERERERERERFVVVURERERERERERDMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzM0RERERERDMzM0RERERERERERGZmZmZmZlVVVVVVVURERFVVVURERERERERERERERERERERERERERERERERERFVVVURERERERERERERERERERFVVVVVVVURERERERERERERERERERFVVVVVVVVVVVVVVVVVVVURERFVVVWZmZlVVVWZmZoiIiIiIiIiIiIiIiHd3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZlVVVURERFVVVVVVVURERERERGZmZmZmZlVVVTMzMzMzMzMzM0RERERERDMzM0RERDMzMzMzM0RERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERGZmZjMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMyIiIiIiIiIiIiIiIkRERDMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzM0RERDMzM0RERDMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMyIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIjMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERERERERERERERDMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIhERESIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIjMzM0RERFVVVXd3d4iIiIiIiJmZmaqqqru7u7u7u8zMzN3d3e7u7u7u7v///+7u7v///////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMzMzMy7u7vMzMzMzMzMzMzd3d3d3d3d3d3u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3u7u7d3d3u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMy7u7u7u7uqqqqqqqqqqqqZmZmZmZmqqqqqqqqqqqqqqqqqqqq7u7u7u7u7u7vMzMzMzMzd3d3MzMzd3d3MzMzd3d3d3d3d3d3MzMzd3d3d3d3MzMzd3d3d3d3MzMzMzMzMzMzMzMzMzMzMzMzd3d3MzMzMzMzMzMzMzMy7u7vMzMzMzMy7u7u7u7u7u7uqqqq7u7u7u7uqqqrMzMzd3d3MzMzMzMzMzMzd3d3d3d3u7u7d3d3d3d3d3d3MzMy7u7uqqqqZmZmqqqqZmZmqqqqqqqqqqqrMzMzMzMzu7u7u7u7u7u7////////////////////////////////////////////u7u7////////////////////////////////////////////u7u7////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7d3d3d3d3d3d3MzMzd3d3u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7d3d3u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3MzMzMzMzd3d3MzMzd3d3MzMzd3d3d3d3d3d3MzMzd3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMy7u7u7u7uqqqqqqqqqqqqqqqqqqqqqqqqqqqqZmZmqqqqZmZmZmZmqqqqZmZmZmZmqqqqqqqqZmZmqqqqZmZmIiIiZmZmIiIiZmZmZmZmIiIiZmZmZmZmZmZmZmZmZmZmZmZmZmZmqqqqIiIiIiIh3d3dmZmZVVVVEREREREREREQzMzNEREREREREREREREQzMzNERERVVVVERERVVVVVVVVERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERVVVVERERERERERERVVVVVVVVVVVVERERVVVVVVVVmZmaIiIiIiIiZmZl3d3dVVVUzMzMzMzMzMzMzMzMiIiIREREREREREREREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMiIiIiIiIREREiIiIzMzMiIiIzMzMzMzMiIiIzMzMzMzNEREQzMzMzMzMiIiIiIiIiIiIzMzMzMzMzMzNEREREREREREQzMzMzMzNEREREREREREQzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNERERmZmZmZmZVVVVEREQzMzNEREREREQzMzMzMzNERERERERERERERERERERERERERERERERVVVVVVVVERERERERERERERERmZmZVVVVEREQzMzMzMzNEREREREQzMzMzMzNERERERERERERERERVVVVEREREREREREQzMzMiIiIiIiIiIiJEREQzMzMiIiIzMzMzMzMiIiIzMzNERERERERERERVVVVERERERERERERERERERERERERERERERERVVVVmZmZmZmZVVVVVVVVERERERERERERVVVVVVVVmZmZVVVVmZmZmZmZmZmZVVVVVVVVERERVVVVEREQzMzMzMzMzMzNERERERERERERVVVVEREREREREREREREREREREREREREREREREREREREREREQzMzMzMzMzMzMzMzNERERERERVVVVEREREREQiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzNEREQzMzMzMzMzMzNERERVVVVVVVVEREREREQzMzMzMzNERERERERVVVVVVVVERERERERERERERERERERVVVVERERVVVVERERVVVVEREREREQzMzMzMzMzMzNVVVVVVVVERERERERVVVVVVVVEREQzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIzMzMzMzMzMzNEREQzMzNEREQzMzMzMzMiIiIzMzNERERERERERERVVVVEREQzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERERERVVVVERERERERERERERERERERERERERERVVVVERERVVVVERERVVVVVVVVERERVVVVVVVVEREREREREREQzMzNEREREREREREREREQzMzNEREQzMzNERERERERVVVVERERERERERERERERERERVVVVmZmZmZmZ3d3dmZmZmZmZVVVVERERERERVVVUzMzNEREREREQzMzNEREQzMzNEREREREQzMzNEREQzMzNEREQzMzMzMzMzMzNEREQzMzMzMzNERERERERVVVVEREQzMzMzMzMzMzNERERERERVVVVmZmZmZmZVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVUzMzMzMzMzMzNERERERERERERERERERERVVVVERERVVVVERERVVVVVVVVEREREREREREREREREREREREREREREREREREQzMzNERERmZmZVVVUzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERVVVVmZmZVVVVERERVVVVVVVVVVVVERERERERERERERERERERERERERERERERERERERERERERVVVVVVVVmZmZVVVVERERERERERERVVVVVVVVERERERERVVVVVVVVVVVVEREQzMzMzMzNERERERERmZmaZmZmZmZmIiIiIiIh3d3d3d3eIiIiIiIh3d3dmZmZmZmZmZmZmZmZVVVVmZmZVVVVERERVVVVERERVVVVmZmZVVVUzMzMzMzNEREQzMzNEREREREQzMzMzMzNEREREREREREREREREREQzMzMzMzNEREREREREREQzMzNERERVVVVEREQzMzMiIiIzMzMiIiIzMzMiIiIzMzMzMzMzMzNEREREREQzMzMiIiIiIiIiIiIzMzMzMzMzMzMzMzNEREQzMzMiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNEREQzMzMzMzMiIiIiIiIzMzMiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMzMzMiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzNERERmZmZ3d3d3d3d3d3eZmZmZmZm7u7vMzMzMzMzd3d3u7u7////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////7u7u////////////////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3dzMzMzMzMzMzMu7u7u7u7zMzMzMzMzMzMzMzMzMzMzMzM3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d7u7u3d3d7u7u3d3d3d3d3d3d3d3dzMzMu7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqmZmZmZmZmZmZqqqqqqqqqqqqu7u7u7u7zMzMzMzMzMzMzMzM3d3d3d3d3d3d3d3dzMzM3d3dzMzMzMzMzMzMzMzMzMzMu7u7zMzMzMzMzMzMu7u7zMzMzMzM3d3d3d3dzMzMzMzMu7u7u7u7u7u7u7u7u7u7u7u7zMzMzMzMu7u7u7u7zMzMzMzMzMzMzMzMzMzM3d3d3d3d3d3dzMzMzMzMzMzMu7u7u7u7mZmZmZmZqqqqqqqqqqqqqqqqu7u7zMzM3d3d7u7u7u7u7u7u7u7u////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u////7u7u////7u7u7u7u7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3d7u7u3d3d7u7u3d3d7u7u3d3d7u7u3d3d7u7u3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzM3d3dzMzMzMzMzMzMu7u7zMzMu7u7zMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7qqqqu7u7u7u7qqqqu7u7qqqqqqqqqqqqmZmZmZmZqqqqmZmZmZmZmZmZiIiIiIiId3d3ZmZmVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmVVVVVVVVZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREREREMzMzREREMzMzMzMzREREREREREREREREREREVVVVREREREREREREVVVVVVVVVVVVMzMzMzMzMzMzREREMzMzIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiERERIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzREREMzMzIiIiMzMzMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVREREMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREVVVVVVVVVVVVVVVVREREREREREREMzMzMzMzMzMzMzMzREREREREREREREREREREREREVVVVVVVVREREMzMzREREREREVVVVREREREREREREMzMzREREREREMzMzMzMzMzMzREREREREVVVVREREREREREREMzMzMzMzIiIiMzMzMzMzREREREREMzMzIiIiMzMzMzMzIiIiMzMzREREMzMzREREVVVVREREVVVVVVVVZmZmZmZmREREREREVVVVVVVVZmZmZmZmVVVVREREREREREREREREVVVVREREVVVVZmZmVVVVVVVVVVVVREREREREREREREREMzMzMzMzREREREREREREVVVVREREREREREREREREREREREREREREVVVVREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVVVVVMzMzIiIiMzMzIiIiMzMzMzMzMzMzREREREREREREMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzREREMzMzREREREREZmZmZmZmVVVVVVVVREREREREVVVVREREREREREREREREREREREREREREVVVVREREVVVVREREVVVVVVVVREREMzMzMzMzIiIiMzMzVVVVVVVVREREREREREREVVVVREREMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREREREREREMzMzIiIiMzMzMzMzREREVVVVREREREREREREMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREREREREREREREREREREREREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREMzMzMzMzREREREREREREREREREREREREREREVVVVVVVVREREMzMzREREVVVVVVVVVVVVZmZmZmZmZmZmVVVVREREVVVVVVVVREREREREREREVVVVREREREREREREREREMzMzREREMzMzREREMzMzREREMzMzMzMzREREMzMzMzMzMzMzREREREREMzMzMzMzMzMzREREREREVVVVVVVVVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVREREVVVVREREVVVVVVVVVVVVVVVVREREREREMzMzMzMzMzMzREREREREREREVVVVVVVVVVVVVVVVVVVVREREREREVVVVREREREREREREREREREREREREREREREREMzMzMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREMzMzREREREREREREREREREREREREREREVVVVREREREREREREREREMzMzREREREREREREVVVVREREREREVVVVd3d3d3d3VVVVREREREREVVVVREREVVVVREREREREREREREREMzMzREREMzMzREREMzMzREREZmZmiIiId3d3ZmZmZmZmZmZmd3d3iIiId3d3d3d3d3d3iIiId3d3ZmZmVVVVREREVVVVVVVVREREVVVVVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREREREREREREREREREREREREREMzMzIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzMzMzIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzREREMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzREREIiIiMzMzIiIiMzMzMzMzMzMzREREVVVVREREMzMzIiIiIiIiIiIiMzMzMzMzIiIiMzMzMzMzMzMzREREMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiREREVVVVVVVVZmZmd3d3iIiImZmZqqqqzMzMzMzM3d3d3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////+7u7u7u7v///+7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3czMzN3d3d3d3d3d3czMzN3d3czMzN3d3e7u7t3d3d3d3czMzMzMzN3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3d3d3czMzN3d3czMzLu7u8zMzLu7u6qqqqqqqqqqqqqqqpmZmaqqqqqqqru7u6qqqqqqqru7u7u7u8zMzMzMzMzMzMzMzMzMzMzMzN3d3czMzMzMzMzMzMzMzMzMzLu7u8zMzLu7u6qqqru7u8zMzN3d3czMzLu7u8zMzMzMzMzMzMzMzLu7u7u7u8zMzLu7u7u7u8zMzMzMzMzMzLu7u7u7u7u7u7u7u8zMzLu7u7u7u8zMzMzMzN3d3d3d3czMzLu7u8zMzMzMzLu7u6qqqqqqqqqqqqqqqpmZmaqqqru7u8zMzMzMzN3d3d3d3e7u7u7u7v///////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7v///+7u7v///+7u7v///+7u7v///+7u7v///////+7u7v///+7u7v///+7u7v///+7u7v///+7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3d3d3e7u7t3d3d3d3d3d3d3d3czMzMzMzN3d3czMzMzMzMzMzMzMzLu7u8zMzLu7u8zMzLu7u8zMzMzMzMzMzMzMzMzMzN3d3czMzMzMzMzMzLu7u7u7u7u7u6qqqoiIiJmZmYiIiHd3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVURERERERFVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d2ZmZmZmZnd3d2ZmZlVVVVVVVURERFVVVURERERERERERERERERERERERFVVVWZmZlVVVURERERERERERERERDMzMzMzMyIiIiIiIiIiIjMzMyIiIjMzMzMzMyIiIhERESIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzM0RERDMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM0RERFVVVTMzM0RERERERERERERERCIiIjMzMzMzM0RERFVVVURERERERERERERERFVVVURERERERGZmZlVVVURERERERERERDMzM0RERERERERERERERFVVVVVVVURERERERERERERERDMzMzMzM0RERERERDMzM0RERERERDMzM0RERERERDMzMzMzMzMzM0RERERERERERERERERERERERERERERERDMzMzMzM0RERERERERERFVVVURERDMzMzMzM0RERDMzM1VVVVVVVVVVVVVVVWZmZnd3d3d3d4iIiJmZmXd3d1VVVURERERERDMzM2ZmZmZmZlVVVURERERERERERFVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVURERFVVVURERERERERERDMzM0RERERERERERFVVVVVVVURERERERDMzM0RERDMzM0RERERERERERERERERERDMzMzMzM0RERDMzMzMzMzMzMyIiIjMzM1VVVVVVVURERDMzMzMzMzMzMzMzMyIiIjMzM0RERERERERERDMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzM1VVVWZmZmZmZlVVVURERERERFVVVURERERERERERERERFVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVURERERERCIiIiIiIiIiIjMzM1VVVVVVVURERFVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERFVVVTMzMzMzMzMzM0RERERERFVVVVVVVURERERERDMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIjMzMzMzM0RERDMzMzMzM0RERERERERERERERERERERERERERFVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVURERDMzMzMzM0RERDMzM0RERERERERERERERFVVVURERERERERERERERERERERERFVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVURERERERERERFVVVURERFVVVURERDMzM0RERDMzM0RERDMzM0RERDMzMzMzM0RERDMzMzMzMzMzM0RERERERERERERERFVVVURERERERERERFVVVVVVVURERFVVVWZmZlVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVURERFVVVVVVVVVVVURERERERERERDMzM0RERERERERERFVVVVVVVVVVVVVVVURERERERFVVVURERFVVVURERERERERERERERERERERERERERDMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzM0RERERERDMzMzMzM0RERERERFVVVURERERERERERFVVVURERDMzMzMzM0RERERERERERERERERERERERERERERERHd3d3d3d1VVVURERERERFVVVURERFVVVWZmZkRERERERDMzM0RERDMzM0RERERERDMzM0RERFVVVWZmZmZmZlVVVURERFVVVVVVVWZmZnd3d2ZmZnd3d4iIiIiIiHd3d2ZmZlVVVURERFVVVURERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERFVVVURERERERERERERERERERDMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMyIiIjMzMzMzM0RERERERDMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERERERERERDMzMzMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzM0RERERERDMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIjMzMyIiIiIiIiIiIjMzM0RERERERDMzMzMzMyIiIjMzMzMzM1VVVVVVVTMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzMyIiIiIiIjMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVXd3d4iIiKqqqqqqqru7u8zMzMzMzO7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7d3d3u7u7u7u7d3d3u7u7u7u7d3d3d3d3d3d3d3d3MzMzd3d3d3d3MzMzMzMzMzMzMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMy7u7u7u7u7u7u7u7uqqqqqqqqqqqqqqqq7u7uqqqq7u7uqqqq7u7u7u7vMzMzMzMzd3d3MzMzd3d3MzMzMzMzMzMy7u7u7u7u7u7u7u7vMzMy7u7u7u7u7u7u7u7vMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMy7u7vMzMy7u7u7u7u7u7u7u7u7u7u7u7u7u7uqqqqqqqq7u7uqqqqqqqq7u7u7u7vMzMzMzMzMzMzMzMy7u7vMzMyqqqqqqqqZmZmZmZmZmZmZmZmZmZmqqqq7u7vMzMzMzMzd3d3u7u7u7u7u7u7////u7u7////u7u7////////////////////////////////////////////////////////////u7u7////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3MzMzMzMzMzMy7u7vMzMzMzMzMzMzMzMzd3d3d3d3d3d3d3d3MzMy7u7u7u7uIiIh3d3dmZmZ3d3dmZmZmZmZmZmZERERVVVVVVVVVVVVVVVVERERVVVVmZmZ3d3dmZmZ3d3d3d3d3d3d3d3dmZmZmZmZmZmZ3d3d3d3d3d3d3d3dmZmZ3d3dmZmZmZmZ3d3dmZmZmZmZVVVVVVVVVVVVVVVVmZmZVVVVERERVVVVVVVVVVVVEREQzMzMzMzMzMzNEREREREQzMzMzMzMiIiIzMzMzMzMiIiIiIiIzMzMiIiIiIiIiIiIiIiIzMzMiIiJEREQzMzMiIiIiIiIzMzNEREQzMzMiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMzMzMiIiIzMzMzMzNEREREREQzMzMzMzMzMzMzMzNEREREREQzMzMzMzMiIiIzMzNEREQzMzNEREREREQzMzNEREQzMzNEREQzMzNEREREREREREREREREREQzMzMzMzMzMzMzMzNERERERERERERERERERERVVVVVVVVERERERERVVVVmZmZVVVVEREQzMzMzMzNERERVVVVERERERERVVVVVVVVERERVVVVERERVVVVEREQzMzNEREQzMzMzMzNEREQzMzNEREREREQzMzMzMzNEREQzMzNERERERERERERERERERERERERERERERERERERERERERERERERVVVVERERERERERERVVVVVVVVmZmZmZmZ3d3dmZmZmZmZVVVVmZmZmZmZ3d3eIiIh3d3dEREQzMzMzMzNERERERERVVVVVVVVVVVVERERERERVVVVVVVVmZmZmZmZVVVVmZmZVVVVVVVVVVVVEREQzMzNERERERERVVVVVVVVERERERERERERERERVVVVEREREREREREREREREREREREREREQzMzNEREQzMzNEREREREQzMzMzMzMiIiIzMzMzMzMzMzNVVVVVVVVEREQzMzMzMzNEREQzMzMzMzNEREREREQzMzMzMzMzMzMiIiIiIiIzMzMzMzNEREQzMzMzMzNEREQzMzNEREQzMzMzMzNERERERERVVVVVVVVVVVVERERERERERERERERVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzNERERmZmZVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREREREQzMzMzMzMzMzMzMzNERERVVVVVVVVEREQzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiJEREREREREREQzMzMzMzNERERERERERERERERVVVVERERERERERERERERVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVEREREREQzMzMzMzNERERERERERERERERERERERERERERVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZVVVVERERVVVVERERVVVVVVVVVVVVEREREREQzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzNERERVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVERERVVVVERERVVVVERERVVVVVVVVmZmZVVVVEREREREQzMzNEREQzMzNERERERERVVVVVVVVERERERERVVVVEREREREREREREREREREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzNEREQzMzMzMzNEREREREREREQzMzMzMzNERERmZmZVVVVVVVVEREREREQzMzMzMzMzMzNERERERERERERERERERERERERERERVVVVmZmZVVVVVVVVVVVVERERVVVVmZmZmZmZEREREREQzMzNERERERERERERERERERERERERERERVVVVVVVVERERERERERERERERVVVVVVVVVVVVmZmZmZmaIiIiZmZmIiIhmZmZVVVVERERVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzNERERERERERERERERVVVVVVVVVVVVEREREREREREQzMzMzMzMzMzMiIiIzMzMzMzNEREQzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIzMzMzMzNERERVVVUzMzMzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzNEREQzMzNEREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNEREREREREREQzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIzMzNVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERmZmZ3d3eIiIiZmZmqqqq7u7vMzMzd3d3d3d3u7u7////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////7u7u3d3dzMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzM3d3dzMzM3d3d3d3d3d3dzMzM3d3dzMzM3d3dzMzM3d3d3d3d3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d7u7u3d3dzMzMzMzMzMzMu7u7u7u7u7u7u7u7qqqqqqqqmZmZqqqqqqqqqqqqqqqqu7u7u7u7zMzMzMzMu7u7zMzMzMzMzMzMzMzMzMzMu7u7qqqqqqqqu7u7u7u7u7u7u7u7zMzMzMzMzMzM3d3d3d3dzMzMzMzMzMzMzMzMu7u7u7u7qqqqu7u7mZmZmZmZmZmZmZmZmZmZiIiIiIiImZmZqqqqu7u7qqqqu7u7zMzMu7u7u7u7u7u7u7u7u7u7qqqqmZmZmZmZmZmZmZmZiIiImZmZmZmZqqqqu7u7zMzMzMzMzMzM3d3dzMzM3d3d3d3d3d3d7u7u7u7u7u7u////////7u7u////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u////3d3d3d3d3d3dzMzMu7u7zMzMzMzMzMzMzMzM3d3dzMzM3d3dzMzMqqqqd3d3VVVVVVVVREREREREVVVVVVVVREREREREREREREREREREVVVVVVVVZmZmZmZmd3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmd3d3d3d3ZmZmd3d3ZmZmd3d3d3d3ZmZmZmZmZmZmVVVVZmZmZmZmiIiImZmZd3d3VVVVVVVVVVVVVVVVREREREREREREREREMzMzMzMzIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiERERIiIiERERIiIiMzMzMzMzREREVVVVREREMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzREREVVVVVVVVREREREREMzMzREREREREMzMzMzMzIiIiMzMzREREREREREREREREREREMzMzREREREREMzMzMzMzREREVVVVREREMzMzMzMzIiIiMzMzREREREREREREREREREREZmZmZmZmZmZmREREREREVVVVREREREREVVVVREREMzMzREREVVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREMzMzMzMzMzMzREREREREMzMzMzMzMzMzREREREREREREREREREREREREREREREREREREREREREREREREREREREREVVVVZmZmZmZmVVVVZmZmVVVVVVVVZmZmVVVVVVVVREREREREREREVVVVREREZmZmVVVVVVVVREREREREREREVVVVZmZmVVVVREREREREVVVVREREVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREVVVVREREREREREREVVVVREREVVVVVVVVREREREREREREREREREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVVVVVVVVVREREREREMzMzMzMzREREMzMzREREMzMzIiIiIiIiMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREMzMzMzMzIiIiMzMzREREVVVVZmZmVVVVVVVVREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVREREREREMzMzMzMzMzMzMzMzVVVVVVVVZmZmVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREMzMzREREREREMzMzIiIiMzMzMzMzMzMzREREREREREREREREREREMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREREREREREVVVVREREREREVVVVVVVVREREVVVVVVVVREREVVVVVVVVVVVVVVVVREREMzMzREREMzMzREREREREREREREREREREREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVMzMzREREMzMzREREREREREREREREREREVVVVREREREREREREVVVVREREVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREMzMzMzMzREREMzMzMzMzREREZmZmZmZmVVVVREREREREMzMzREREREREREREREREREREREREREREREREREREREREVVVVVVVVZmZmREREVVVVVVVVd3d3VVVVREREREREREREREREREREREREREREREREREREREREVVVVREREREREREREVVVVREREREREVVVVVVVVVVVVVVVVZmZmiIiIiIiIiIiIZmZmREREVVVVREREREREREREREREZmZmVVVVREREMzMzMzMzREREMzMzREREREREMzMzREREREREVVVVREREVVVVVVVVVVVVREREMzMzREREREREIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREIiIiMzMzREREMzMzREREMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzIiIiREREREREMzMzMzMzMzMzMzMzMzMzREREMzMzREREVVVVVVVVVVVVVVVVMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREVVVVZmZmiIiImZmZqqqqzMzMzMzM3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////+7u7szMzLu7u7u7u6qqqru7u7u7u7u7u7u7u7u7u7u7u8zMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3e7u7t3d3d3d3e7u7t3d3e7u7u7u7u7u7u7u7t3d3e7u7t3d3e7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3czMzMzMzN3d3czMzMzMzMzMzMzMzMzMzN3d3czMzN3d3czMzN3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3e7u7u7u7u7u7t3d3d3d3czMzMzMzLu7u7u7u6qqqqqqqqqqqpmZmaqqqpmZmaqqqqqqqqqqqqqqqqqqqru7u7u7u7u7u7u7u7u7u6qqqru7u7u7u7u7u7u7u6qqqru7u7u7u7u7u7u7u7u7u7u7u8zMzMzMzMzMzMzMzLu7u7u7u7u7u6qqqpmZmZmZmZmZmZmZmYiIiIiIiIiIiIiIiJmZmZmZmaqqqqqqqru7u7u7u7u7u8zMzLu7u7u7u7u7u7u7u7u7u7u7u5mZmZmZmYiIiIiIiIiIiIiIiJmZmZmZmZmZmYiIiJmZmZmZmZmZmZmZmaqqqqqqqru7u8zMzN3d3d3d3e7u7u7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7t3d3bu7u6qqqru7u7u7u8zMzLu7u8zMzMzMzMzMzKqqqnd3d0RERERERERERERERERERERERERERERERDMzM0RERERERERERERERFVVVWZmZmZmZnd3d4iIiIiIiHd3d3d3d2ZmZmZmZnd3d3d3d2ZmZmZmZmZmZoiIiIiIiIiIiHd3d2ZmZmZmZmZmZnd3d3d3d3d3d2ZmZmZmZlVVVVVVVWZmZmZmZmZmZmZmZlVVVTMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMyIiIiIiIhERESIiIiIiIiIiIjMzM0RERDMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzM1VVVURERERERDMzMzMzM0RERFVVVVVVVURERERERERERDMzMzMzMzMzM0RERERERERERERERERERERERFVVVVVVVURERDMzMyIiIkRERERERERERERERDMzMzMzM0RERDMzM0RERDMzM0RERERERFVVVVVVVWZmZlVVVVVVVURERERERFVVVURERERERDMzM0RERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERDMzM1VVVURERERERERERERERERERDMzM0RERERERFVVVVVVVWZmZlVVVWZmZmZmZmZmZlVVVVVVVURERERERFVVVXd3d3d3d1VVVURERERERERERERERERERFVVVURERERERERERDMzM0RERDMzM0RERGZmZmZmZlVVVURERFVVVWZmZlVVVURERERERFVVVURERFVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERDMzMzMzMzMzM0RERFVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIkRERFVVVWZmZlVVVVVVVURERFVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERDMzM0RERDMzM0RERDMzMzMzMyIiIiIiIjMzM0RERFVVVVVVVVVVVURERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVURERDMzMzMzMzMzMzMzM0RERFVVVVVVVURERERERERERDMzMzMzMzMzM0RERDMzM0RERERERERERDMzMzMzM0RERDMzM0RERDMzMyIiIjMzM0RERDMzM0RERERERERERFVVVURERDMzMzMzM0RERERERERERDMzMyIiIjMzMzMzMzMzMyIiIiIiIjMzMyIiIiIiIjMzMzMzM0RERERERERERERERDMzM0RERERERERERERERFVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERDMzM0RERDMzM0RERERERERERERERFVVVURERFVVVURERERERERERFVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERGZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVURERFVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZnd3d3d3d2ZmZmZmZlVVVVVVVVVVVVVVVWZmZlVVVVVVVWZmZlVVVVVVVVVVVTMzMzMzM0RERERERERERERERFVVVVVVVVVVVVVVVURERERERFVVVVVVVURERFVVVVVVVURERERERERERDMzMyIiIjMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMyIiIjMzMzMzMzMzMzMzMyIiIiIiIkRERFVVVVVVVURERDMzM0RERDMzM0RERDMzM0RERERERERERERERERERERERERERERERFVVVWZmZlVVVVVVVVVVVWZmZkRERERERERERERERERERDMzMzMzM0RERERERFVVVVVVVURERDMzM0RERERERERERERERFVVVWZmZmZmZkRERDMzM0RERERERFVVVWZmZmZmZmZmZmZmZnd3d3d3d3d3d0RERFVVVWZmZkRERDMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERERERDMzMzMzMzMzM0RERERERDMzMyIiIiIiIjMzMzMzM0RERFVVVTMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzMzMzM0RERDMzM0RERERERFVVVURERDMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzM0RERERERFVVVTMzMzMzMyIiIjMzMyIiIjMzMzMzMyIiIjMzMyIiIjMzMyIiIiIiIjMzMyIiIiIiIjMzM0RERDMzM0RERERERERERERERFVVVVVVVVVVVURERDMzMzMzMzMzM0RERDMzMyIiIiIiIiIiIjMzMyIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERFVVVWZmZnd3d4iIiJmZmbu7u8zMzMzMzN3d3e7u7v///+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////u7u7d3d3MzMzMzMzMzMy7u7u7u7u7u7u7u7uZmZmZmZmZmZmqqqqqqqqqqqq7u7u7u7vMzMzMzMzMzMzd3d3MzMzd3d3d3d3d3d3d3d3u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7d3d3d3d3u7u7d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMzMzMzd3d3MzMzMzMzd3d3d3d3d3d3d3d3MzMzd3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMy7u7u7u7uqqqqqqqqqqqqqqqqqqqq7u7uqqqqqqqqZmZmZmZmqqqqqqqq7u7uqqqq7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7uqqqq7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7uqqqqqqqqqqqqZmZmIiIiIiIiIiIiIiIiZmZmqqqqqqqqqqqqqqqqqqqqqqqq7u7u7u7u7u7u7u7u7u7vMzMy7u7u7u7u7u7u7u7uqqqqqqqqqqqqZmZmIiIiIiIiIiIh3d3eIiIiIiIiZmZmIiIiIiIiIiIh3d3eIiIiIiIiqqqqqqqq7u7vMzMzd3d3d3d3u7u7u7u7u7u7////u7u7////////////////////////////////////////////////////////////////////////////////////////u7u7////////u7u7////////////u7u7////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////u7u7////////////u7u7////u7u7////////u7u7u7u7u7u7d3d3MzMzMzMyqqqq7u7vMzMzMzMzMzMzMzMzd3d3MzMy7u7uZmZlVVVVVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNERERVVVVVVVVmZmZ3d3eIiIh3d3d3d3dmZmZmZmZmZmZ3d3dmZmZmZmZVVVVmZmZ3d3eZmZl3d3dmZmZVVVVVVVVmZmZmZmZVVVVEREQzMzNERERERERVVVVmZmZ3d3eZmZl3d3dVVVUzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIzMzMzMzMiIiIzMzNEREQzMzMzMzMzMzMzMzNERERVVVVEREREREQzMzMzMzNERERERERERERERERERERVVVVVVVVVVVVVVVVEREREREQzMzMzMzMzMzNERERVVVVEREREREQzMzNEREQzMzMzMzNERERERERVVVVVVVVVVVVVVVVVVVVmZmZEREREREREREREREQzMzNEREQzMzNERERVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVERERVVVVERERmZmZmZmZVVVVERERERERERERVVVVVVVVVVVVVVVVmZmZ3d3d3d3d3d3d3d3d3d3dmZmZVVVVERERERERERERVVVV3d3dVVVVERERERERERERERERVVVVVVVVVVVVEREREREREREREREQzMzNERERERERmZmZ3d3d3d3dVVVVmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVERERVVVVVVVVEREREREREREREREREREREREQzMzMzMzMzMzNERERVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVEREREREREREQzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERmZmZmZmZVVVVmZmZVVVVEREREREREREQzMzMzMzMzMzNEREQzMzNEREQzMzNEREQzMzMzMzNEREQzMzMzMzMiIiIzMzMzMzNERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVVEREREREQzMzMzMzMzMzNERERVVVVERERERERVVVVVVVVEREQzMzMzMzMzMzMzMzNEREREREREREQzMzNEREQzMzMzMzNEREQzMzMiIiIzMzNEREQzMzMzMzNERERERERERERVVVVEREQzMzMzMzNEREREREQzMzMzMzMzMzNEREREREQzMzMzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzNEREQzMzNERERERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVEREQzMzNEREQzMzMzMzNEREREREQzMzMzMzNERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVEREQzMzMzMzMzMzMzMzNEREREREQzMzNERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZ3d3d3d3d3d3d3d3dVVVVVVVVmZmZVVVVmZmZmZmZVVVVVVVVmZmZVVVVERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVERERERERVVVVERERVVVVVVVVVVVVmZmZEREREREQzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzNERERVVVVERERERERERERERERERERERERERERERERERERERERERERVVVVVVVVVVVVERERVVVVmZmZmZmZVVVVVVVVEREREREREREREREREREQzMzNEREQzMzNEREREREREREREREREREQzMzMzMzNERERVVVVEREREREREREQzMzMzMzMzMzNEREQzMzNERERVVVVVVVV3d3eIiIiqqqp3d3czMzNEREREREQzMzNEREQzMzMzMzMzMzMzMzNEREREREREREREREREREREREQzMzMzMzMiIiIzMzNEREREREREREREREQzMzMzMzMzMzMzMzNEREREREREREQzMzMzMzNEREQzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREQzMzNEREREREREREREREQiIiIzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIzMzMiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzNEREREREREREREREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVEREREREREREREREQzMzMzMzMiIiIzMzMiIiIiIiJERERERERERERVVVV3d3d3d3eIiIiIiIiqqqq7u7vMzMzMzMzd3d3u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////7u7u7u7u7u7u7u7u3d3d7u7u3d3d7u7u3d3d3d3dzMzMzMzMu7u7u7u7qqqqqqqqu7u7u7u7qqqqqqqqqqqqu7u7u7u7u7u7u7u7zMzMu7u7zMzMzMzMzMzM3d3d3d3d7u7u7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzM3d3dzMzMzMzMzMzM3d3dzMzM3d3d3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMu7u7qqqqu7u7u7u7qqqqu7u7qqqqmZmZmZmZmZmZmZmZmZmZqqqqqqqqqqqqu7u7qqqqzMzMzMzMu7u7u7u7u7u7u7u7qqqqqqqqu7u7qqqqqqqqqqqqu7u7qqqqqqqqqqqqqqqqqqqqmZmZmZmZmZmZmZmZqqqqqqqqu7u7u7u7qqqqqqqqqqqqqqqqqqqqqqqqu7u7u7u7zMzMu7u7zMzMzMzMzMzMu7u7qqqqqqqqqqqqqqqqiIiId3d3iIiIiIiIiIiIiIiIiIiId3d3ZmZmZmZmZmZmZmZmZmZmd3d3d3d3iIiIiIiIqqqqu7u7zMzM3d3d7u7u////7u7u////////////7u7u////////7u7u////////////7u7u////////////////////7u7u////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////7u7u////////////7u7u////////////////////////////////////////////////////////7u7u////////////////////////////////////////////7u7u////7u7u////7u7u7u7u7u7u7u7u3d3dzMzM3d3dzMzMzMzMu7u7qqqqqqqqu7u7u7u7u7u7zMzM3d3d3d3d3d3d3d3dzMzMmZmZd3d3VVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzREREREREVVVVVVVVZmZmZmZmZmZmVVVVZmZmVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVZmZmVVVVVVVVREREMzMzMzMzREREREREVVVVVVVVZmZmiIiIZmZmVVVVMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiERERIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiREREREREREREMzMzIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREREREMzMzIiIiMzMzMzMzVVVVMzMzMzMzREREMzMzREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVREREREREMzMzREREREREVVVVVVVVVVVVREREREREMzMzMzMzREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVREREREREVVVVREREREREREREREREREREVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmVVVVREREREREd3d3iIiIZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmVVVVZmZmZmZmVVVVREREMzMzMzMzREREZmZmVVVVREREREREVVVVVVVVREREREREVVVVVVVVREREREREMzMzREREREREREREVVVVZmZmd3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREREREREREREREVVVVVVVVVVVVREREREREREREREREREREREREREREREREMzMzMzMzREREVVVVZmZmZmZmZmZmVVVVVVVVVVVVREREREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzMzMzMzMzMzMzREREVVVVVVVVVVVVREREREREMzMzMzMzMzMzREREREREREREREREREREREREMzMzMzMzREREMzMzMzMzMzMzMzMzIiIiMzMzREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREMzMzMzMzMzMzREREVVVVREREREREVVVVVVVVREREVVVVREREREREMzMzREREREREVVVVVVVVREREREREMzMzMzMzREREMzMzMzMzMzMzREREREREMzMzREREREREREREMzMzMzMzMzMzREREREREREREREREREREVVVVREREMzMzREREMzMzMzMzMzMzIiIiMzMzREREREREMzMzREREREREREREREREVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVREREREREMzMzMzMzMzMzMzMzMzMzREREREREREREREREVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVREREVVVVZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmREREREREMzMzMzMzMzMzMzMzREREREREMzMzREREREREREREMzMzMzMzREREREREVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmVVVVZmZmVVVVVVVVVVVVMzMzREREREREREREREREVVVVVVVVZmZmZmZmVVVVREREREREREREREREVVVVVVVVVVVVVVVVVVVVREREREREREREMzMzIiIiREREREREREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREMzMzMzMzREREMzMzMzMzREREMzMzMzMzREREREREVVVVREREREREREREREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVREREZmZmZmZmREREVVVVREREREREMzMzREREREREREREMzMzMzMzREREREREREREMzMzREREREREVVVVZmZmVVVVREREMzMzIiIiIiIiMzMzIiIiMzMzMzMzREREMzMzZmZmqqqqqqqqZmZmMzMzREREMzMzMzMzREREMzMzREREREREREREREREVVVVREREREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREVVVVVVVVREREREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiMzMzMzMzIiIiIiIiREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzIiIiMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzMzMzREREMzMzREREREREREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREREREMzMzMzMzIiIiMzMzIiIiIiIiIiIiMzMzMzMzIiIiMzMzMzMzIiIiIiIiIiIiMzMzIiIiIiIiMzMzIiIiIiIiMzMzIiIiMzMzREREREREREREVVVVVVVVVVVVVVVVREREMzMzMzMzMwD//wAAMzMzMzMiIiIzMzNERERERERVVVVmZmZ3d3eIiIiZmZmqqqqqqqrMzMzMzMzd3d3u7u7u7u7////////u7u7////////u7u7////////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u7u7u3d3d3d3d3d3d3d3du7u7zMzMzMzMu7u7zMzMu7u7zMzMu7u7zMzMzMzM3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzM3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM3d3dzMzMzMzM3d3d3d3d3d3dzMzMzMzM3d3dzMzM3d3d3d3dzMzMzMzMzMzMzMzMu7u7u7u7u7u7qqqqqqqqmZmZmZmZqqqqmZmZmZmZqqqqmZmZqqqqqqqqqqqqqqqqu7u7qqqqu7u7qqqqqqqqqqqqqqqqmZmZmZmZiIiImZmZmZmZqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqu7u7u7u7qqqqqqqqqqqqmZmZmZmZqqqqu7u7qqqqqqqqu7u7u7u7u7u7u7u7u7u7zMzMu7u7qqqqqqqqmZmZmZmZiIiIiIiIiIiIiIiId3d3d3d3ZmZmVVVVVVVVVVVVVVVVREREREREREREREREVVVVZmZmd3d3mZmZqqqqu7u7zMzM3d3d7u7u7u7u////7u7u////////////////////////////7u7u////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3dzMzMzMzMzMzMu7u7u7u7qqqqqqqqu7u7u7u7qqqqu7u7qqqqu7u7u7u7u7u7u7u7zMzMzMzM3d3dzMzMzMzMiIiIZmZmREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmVVVVREREREREREREREREREREREREREREREREMzMzREREMzMzMzMzREREREREMzMzIiIiMzMzMzMzIiIiERERIiIiMzMzIiIiIiIiIiIiIiIiIiIiERERERERERERIiIiIiIiIiIiIiIiREREZmZmZmZmVVVVREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREMzMzREREREREVVVVVVVVVVVVZmZmZmZmZmZmREREREREREREVVVVVVVVREREREREREREREREREREREREREREREREREREVVVVVVVVZmZmZmZmZmZmVVVVVVVVREREVVVVREREREREREREVVVVVVVVVVVVZmZmiIiIiIiIiIiIiIiImZmZqqqqd3d3VVVVVVVVVVVVVVVVd3d3iIiId3d3ZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVZmZmREREMzMzMzMzREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVREREMzMzMzMzMzMzMzMzVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREREREREREREREREREREREREREREREVVVVZmZmd3d3ZmZmVVVVREREREREVVVVVVVVREREMzMzMzMzMzMzIiIiMzMzREREREREREREREREREREMzMzREREMzMzIiIiIiIiMzMzREREREREREREREREMzMzMzMzMzMzREREREREREREMzMzREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzVVVVVVVVVVVVVVVVREREVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmVVVVREREVVVVVVVVREREREREREREREREVVVVREREREREREREVVVVZmZmVVVVREREVVVVREREREREVVVVVVVVVVVVREREREREMzMzREREREREMzMzREREREREREREREREREREREREREREMzMzREREREREVVVVREREREREREREREREVVVVREREREREMzMzREREREREMzMzMzMzMzMzVVVVVVVVREREREREREREREREVVVVVVVVVVVVd3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVREREREREREREREREREREREREREREREREREREREREVVVVREREREREVVVVVVVVZmZmVVVVREREVVVVREREVVVVVVVVVVVVREREVVVVREREREREZmZmVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREREREMzMzREREVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVZmZmVVVVZmZmVVVVVVVVZmZmVVVVVVVVREREREREREREVVVVREREREREVVVVVVVVREREVVVVREREMzMzREREREREREREREREREREVVVVREREREREREREREREMzMzMzMzIiIiREREREREMzMzREREREREREREREREMzMzMzMzREREMzMzREREREREMzMzREREMzMzREREREREVVVVREREREREIiIiMzMzVVVVVVVVVVVVREREREREREREREREREREVVVVREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVREREVVVVVVVVREREVVVVREREREREREREMzMzREREMzMzMzMzREREREREMzMzREREREREREREREREZmZmd3d3d3d3VVVVIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzZmZmiIiId3d3VVVVMzMzREREMzMzREREREREREREREREREREVVVVREREREREREREREREREREMzMzMzMzMzMzMzMzREREMzMzREREREREVVVVVVVVZmZmVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiREREMzMzMzMzMzMzMzMzIiIiIiIiMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzMzMzMzMzIiIiMzMzMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiMzMzMzMzIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREVVVVREREVVVVVVVVVVVVREREREREMzMzMzMzIiIiMzMzREREREREVVVVd3d3d3d3iIiImZmZqqqqu7u7u7u7zMzM3d3d7u7u////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////+7u7t3d3e7u7u7u7t3d3d3d3d3d3e7u7t3d3d3d3d3d3e7u7t3d3d3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3d3d3czMzMzMzKqqqru7u7u7u7u7u7u7u7u7u7u7u8zMzN3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzN3d3czMzN3d3czMzMzMzN3d3czMzN3d3d3d3d3d3d3d3czMzMzMzMzMzLu7u7u7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqpmZmaqqqqqqqpmZmaqqqqqqqqqqqqqqqpmZmaqqqpmZmYiIiIiIiJmZmYiIiJmZmYiIiJmZmZmZmaqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqpmZmZmZmaqqqqqqqpmZmaqqqqqqqqqqqpmZmaqqqqqqqqqqqru7u7u7u6qqqru7u6qqqqqqqpmZmaqqqpmZmZmZmYiIiHd3d2ZmZmZmZlVVVVVVVVVVVVVVVURERERERDMzMzMzM0RERERERFVVVWZmZnd3d4iIiJmZmbu7u7u7u93d3d3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////+7u7v///////////+7u7v///+7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3d3d3e7u7t3d3d3d3e7u7t3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzLu7u8zMzLu7u8zMzLu7u8zMzLu7u8zMzMzMzMzMzMzMzMzMzLu7u8zMzLu7u8zMzLu7u7u7u6qqqoiIiFVVVVVVVURERFVVVVVVVWZmZmZmZlVVVVVVVVVVVWZmZlVVVWZmZlVVVURERFVVVWZmZlVVVWZmZlVVVWZmZmZmZnd3d3d3d2ZmZnd3d3d3d2ZmZmZmZnd3d3d3d3d3d3d3d4iIiGZmZlVVVVVVVURERGZmZnd3d1VVVURERERERDMzM0RERDMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERCIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMxERESIiIiIiIhERESIiIhERESIiIhERERERESIiIiIiIiIiIkRERERERGZmZmZmZkRERDMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERDMzM0RERERERERERFVVVVVVVWZmZlVVVXd3d3d3d1VVVURERERERFVVVVVVVVVVVURERERERDMzM0RERERERERERERERERERERERERERFVVVVVVVVVVVWZmZmZmZmZmZlVVVURERERERFVVVVVVVWZmZnd3d3d3d3d3d5mZmYiIiHd3d3d3d4iIiGZmZlVVVURERDMzM1VVVXd3d3d3d1VVVVVVVURERFVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVURERERERERERERERERERERERFVVVWZmZlVVVVVVVWZmZmZmZlVVVWZmZmZmZnd3d1VVVURERFVVVTMzMzMzMzMzM0RERDMzM0RERGZmZmZmZmZmZmZmZmZmZnd3d3d3d1VVVVVVVVVVVVVVVURERERERFVVVURERFVVVURERERERERERERERERERERERFVVVURERFVVVURERFVVVWZmZmZmZlVVVVVVVURERFVVVVVVVURERDMzMzMzMyIiIjMzMzMzM0RERDMzM0RERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVURERDMzMzMzM0RERDMzMzMzMzMzM0RERDMzMzMzM0RERERERERERFVVVURERERERDMzMzMzM0RERERERFVVVURERFVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZlVVVURERFVVVURERFVVVURERERERERERFVVVVVVVVVVVURERFVVVVVVVURERERERERERERERERERERERDMzM0RERERERERERERERERERDMzM0RERERERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVURERERERERERDMzMzMzM0RERDMzMzMzM0RERERERFVVVURERERERERERFVVVVVVVWZmZlVVVVVVVVVVVWZmZmZmZlVVVVVVVWZmZlVVVVVVVVVVVWZmZmZmZlVVVURERFVVVVVVVTMzM0RERERERERERERERERERFVVVURERERERERERFVVVVVVVVVVVVVVVURERERERERERFVVVURERERERFVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVTMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVURERERERFVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZlVVVVVVVURERERERGZmZlVVVURERFVVVVVVVVVVVURERDMzM0RERERERERERERERERERFVVVVVVVURERERERERERERERDMzMzMzMyIiIjMzMzMzMzMzM0RERERERERERDMzMzMzMzMzMzMzM0RERDMzM0RERDMzM0RERDMzM0RERERERERERERERERERCIiIjMzM2ZmZnd3d1VVVVVVVURERERERERERERERERERERERFVVVURERFVVVURERFVVVVVVVVVVVURERERERERERERERFVVVURERFVVVURERERERERERDMzM0RERERERERERERERERERDMzM0RERDMzM1VVVWZmZnd3d2ZmZkRERCIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzM0RERGZmZnd3d1VVVURERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVTMzM0RERERERDMzMzMzMyIiIkRERGZmZlVVVURERDMzM1VVVURERFVVVURERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVTMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIhERERERESIiIhERESIiIjMzMzMzMyIiIjMzM0RERERERERERERERDMzM0RERDMzM0RERERERERERDMzMzMzM0RERERERDMzM0RERERERERERFVVVVVVVVVVVURERERERDMzMzMzMzMzM0RERERERERERFVVVVVVVWZmZnd3d4iIiKqqqru7u8zMzMzMzN3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3MzMzMzMy7u7vMzMy7u7uqqqqqqqqqqqqqqqq7u7u7u7vMzMzMzMzMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3MzMzMzMzMzMzMzMzMzMzMzMzd3d3MzMzMzMzMzMy7u7vMzMzMzMzMzMzd3d3MzMzd3d3MzMzMzMzd3d3d3d3MzMzd3d3MzMzd3d3d3d3MzMzMzMy7u7u7u7u7u7uqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqZmZmZmZmZmZmZmZmIiIiIiIiZmZmZmZmIiIiIiIiIiIiIiIiIiIiZmZmZmZmZmZmqqqqqqqqqqqqqqqqqqqqZmZmqqqqZmZmZmZmZmZmZmZmZmZmZmZmZmZmIiIiIiIiIiIiZmZmZmZmZmZmqqqqqqqq7u7u7u7uqqqq7u7u7u7u7u7uqqqqZmZmIiIiZmZmIiIh3d3dmZmZmZmZVVVVEREREREQzMzMzMzNEREQzMzNERERVVVVVVVVVVVVmZmZ3d3eIiIiZmZmZmZmqqqrMzMzMzMzd3d3u7u7////////////////////u7u7////////////////////////////////////////////////////////////////////////////u7u7////////////u7u7////u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7d3d3u7u7d3d3u7u7d3d3d3d3u7u7d3d3u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3MzMzd3d3d3d3MzMzd3d3MzMzd3d3d3d3d3d3d3d3d3d3MzMzd3d3MzMzd3d3MzMzMzMzMzMy7u7uqqqqqqqqZmZmZmZmIiIh3d3d3d3dVVVVmZmZmZmZ3d3d3d3dmZmZ3d3d3d3dmZmZ3d3d3d3dVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3dmZmZVVVVmZmZmZmZ3d3eIiIiIiIiIiIh3d3dmZmZVVVVERERVVVVVVVVVVVVERERVVVVEREQzMzNEREQzMzMzMzMzMzMiIiIzMzNEREQzMzMzMzMzMzMzMzMzMzMiIiIREREiIiIiIiIzMzMzMzMREREiIiIiIiIiIiIREREiIiIREREREREREREiIiIiIiIREREREREiIiIiIiIzMzNERERVVVVEREQzMzMzMzNEREQzMzNEREQzMzNEREREREQzMzMzMzMzMzNEREQzMzMzMzMzMzNERERERERERERERERERERERERERERERERERERVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVEREQzMzMzMzNVVVV3d3dmZmZVVVVERERVVVVVVVVVVVVmZmZmZmZmZmZVVVV3d3dmZmZVVVVERERVVVV3d3d3d3dmZmZVVVV3d3dmZmZ3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3dmZmZVVVVEREQzMzMiIiJERER3d3dmZmZVVVVVVVVERERVVVVVVVVERERVVVVmZmZmZmZmZmZmZmZVVVVEREQzMzNEREQzMzNERERVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZVVVVEREREREREREQzMzMzMzNEREQzMzNERERVVVVVVVVmZmZmZmZ3d3d3d3d3d3dmZmZVVVVmZmZVVVVVVVVVVVVERERERERVVVVERERERERVVVVVVVVVVVVERERVVVVVVVVVVVVERERERERERERmZmZ3d3dmZmZVVVVVVVVEREREREQzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzNEREREREREREREREQzMzMzMzMzMzNEREQzMzNEREREREQzMzMzMzMzMzNERERVVVVEREREREQzMzMzMzNERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZ3d3dmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZERERERERERERERERERERVVVVVVVVVVVVERERVVVVERERVVVVERERERERVVVVVVVVEREREREQzMzNEREQzMzNERERERERERERERERERERERERERERVVVVVVVVVVVVVVVVERERERERVVVVVVVVERERVVVVEREREREQzMzMzMzMzMzMzMzMzMzNERERVVVVERERERERERERmZmZ3d3dmZmZVVVVVVVVmZmZmZmZ3d3dmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVERERERERERERERERERERVVVVVVVVERERERERVVVVVVVVVVVVmZmZERERVVVVERERERERVVVVERERERERVVVVERERVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVV3d3dmZmZEREQzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVmZmZVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERVVVVVVVVERERERERERERVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREREREQzMzMzMzMzMzMzMzNEREQzMzMzMzNEREQzMzNEREQzMzNEREQzMzMzMzMzMzMzMzNmZmZ3d3dmZmZVVVVERERERERERERERERERERERERVVVVERERVVVVERERVVVVVVVVERERVVVVVVVVERERERERERERERERERERVVVVEREQzMzNEREREREQzMzNERERERERVVVVEREQzMzNERERVVVVmZmZmZmZVVVUzMzMiIiIiIiIzMzMzMzMzMzMzMzNERERVVVVERERVVVVmZmZVVVVERERERERERERERERVVVVVVVVmZmZVVVVVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzNERER3d3dmZmZERERERERVVVVVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNEREREREQzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIREREREREiIiIREREiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzNERERERERERERVVVVEREREREREREREREREREREREREREREREREREREREREREQzMzMzMzNERERERERVVVVVVVVmZmZmZmZEREQzMzMzMzNVVVVERERERERVVVVmZmZVVVVmZmaIiIiqqqqqqqrMzMzMzMzMzMzd3d3u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////7u7u3d3d7u7u7u7u7u7u7u7u3d3d7u7u7u7u3d3d7u7u3d3d3d3d7u7u3d3d3d3d7u7u3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3dzMzMu7u7u7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqqqqqu7u7qqqqu7u7u7u7zMzMu7u7zMzMzMzMzMzM3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzM3d3dzMzM3d3dzMzMzMzM3d3dzMzMzMzMzMzMzMzMzMzMu7u7zMzMu7u7zMzMzMzMzMzMzMzMzMzMzMzM3d3dzMzM3d3dzMzM3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMu7u7u7u7u7u7qqqqqqqqqqqqqqqqu7u7qqqqqqqqqqqqqqqqmZmZmZmZiIiIiIiIiIiIiIiImZmZiIiImZmZiIiImZmZmZmZiIiImZmZmZmZmZmZqqqqqqqqmZmZqqqqqqqqqqqqqqqqmZmZiIiIiIiId3d3d3d3ZmZmd3d3ZmZmZmZmd3d3iIiImZmZmZmZqqqqqqqqqqqqu7u7u7u7qqqqqqqqqqqqqqqqqqqqiIiIiIiIiIiId3d3ZmZmVVVVREREREREMzMzMzMzREREMzMzMzMzREREREREREREZmZmZmZmd3d3ZmZmd3d3d3d3mZmZqqqqu7u7zMzMzMzM3d3d7u7u7u7u////////////////////////////////7u7u////////////////7u7u////7u7u////7u7u7u7u////7u7u////7u7u////7u7u7u7u7u7u7u7u3d3d7u7u3d3d7u7u7u7u7u7u3d3d3d3d3d3d7u7u3d3d7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u7u7u3d3d7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMu7u7u7u7qqqqqqqqiIiImZmZiIiIiIiIZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmVVVVVVVVZmZmREREREREREREREREVVVVREREREREVVVVVVVVREREVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmd3d3d3d3VVVVREREZmZmZmZmVVVVREREREREZmZmiIiIZmZmREREMzMzMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiERERIiIiIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzREREMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREREREREREREREREREREREMzMzMzMzREREREREREREVVVVREREREREREREREREREREZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVMzMzMzMzREREVVVVd3d3iIiId3d3VVVVZmZmZmZmd3d3iIiIiIiIiIiId3d3iIiId3d3ZmZmREREMzMzVVVVd3d3ZmZmZmZmZmZmZmZmZmZmiIiId3d3d3d3d3d3iIiIiIiId3d3d3d3ZmZmMzMzMzMzMzMzVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREMzMzVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVZmZmREREREREREREREREREREREREREREREREREREREREREREVVVVZmZmZmZmd3d3iIiIiIiId3d3ZmZmZmZmd3d3VVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREVVVVZmZmZmZmZmZmVVVVREREREREMzMzMzMzIiIiMzMzREREMzMzREREVVVVVVVVREREREREMzMzMzMzIiIiMzMzMzMzREREREREREREREREMzMzREREMzMzMzMzREREREREREREREREREREREREVVVVVVVVVVVVREREREREREREMzMzREREREREVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmd3d3ZmZmd3d3d3d3d3d3ZmZmVVVVVVVVVVVVVVVVZmZmZmZmREREVVVVREREVVVVREREREREREREREREVVVVVVVVVVVVREREREREREREREREREREREREREREMzMzMzMzREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREREREMzMzREREREREREREMzMzMzMzVVVVVVVVREREREREVVVVZmZmd3d3ZmZmZmZmVVVVZmZmZmZmd3d3ZmZmZmZmVVVVVVVVREREREREVVVVZmZmVVVVVVVVVVVVREREREREVVVVREREREREVVVVREREREREREREREREREREREREVVVVZmZmVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREVVVVZmZmVVVVREREREREMzMzMzMzMzMzREREMzMzREREMzMzREREMzMzVVVVd3d3VVVVZmZmZmZmd3d3ZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVZmZmVVVVVVVVVVVVREREVVVVREREVVVVREREVVVVVVVVVVVVREREREREREREMzMzMzMzMzMzIiIiMzMzMzMzREREVVVVVVVVVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREREREREREZmZmZmZmZmZmVVVVREREREREREREREREREREREREREREREREREREVVVVREREVVVVREREVVVVREREREREREREREREREREREREREREREREREREREREREREREREREREVVVVREREREREMzMzREREREREREREMzMzMzMzMzMzIiIiMzMzMzMzREREREREVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREVVVVVVVVZmZmZmZmVVVVREREMzMzMzMzMzMzMzMzMzMzREREMzMzREREd3d3ZmZmREREVVVVVVVVREREMzMzMzMzMzMzIiIiMzMzMzMzIiIiREREMzMzIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzREREREREREREMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiIiIiIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzREREREREMzMzMzMzMzMzMzMzREREREREVVVVVVVVREREREREMzMzMzMzMzMzREREREREREREVVVVZmZmd3d3ZmZmVVVVREREVVVVREREVVVVVVVVZmZmVVVVZmZmd3d3mZmZqqqqu7u7zMzMzMzMzMzM7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////+7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7t3d3d3d3czMzMzMzO7u7t3d3d3d3d3d3czMzMzMzMzMzLu7u7u7u6qqqqqqqru7u6qqqqqqqqqqqqqqqqqqqpmZmaqqqqqqqqqqqru7u6qqqru7u7u7u8zMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzN3d3czMzMzMzMzMzN3d3czMzMzMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u7u7u8zMzMzMzMzMzN3d3czMzMzMzN3d3d3d3czMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u6qqqru7u6qqqru7u7u7u7u7u7u7u6qqqqqqqpmZmYiIiIiIiIiIiIiIiJmZmZmZmZmZmYiIiIiIiIiIiJmZmYiIiIiIiJmZmYiIiIiIiJmZmaqqqpmZmaqqqpmZmYiIiHd3d3d3d3d3d2ZmZmZmZmZmZmZmZoiIiHd3d4iIiIiIiIiIiJmZmZmZmZmZmaqqqqqqqqqqqqqqqpmZmaqqqpmZmaqqqpmZmYiIiHd3d3d3d2ZmZlVVVURERERERERERERERERERERERERERDMzM0RERFVVVURERERERFVVVURERFVVVURERFVVVWZmZnd3d5mZmbu7u8zMzN3d3e7u7u7u7v///+7u7v///+7u7v///+7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3e7u7u7u7t3d3e7u7t3d3d3d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzLu7u7u7u6qqqpmZmZmZmYiIiHd3d2ZmZlVVVVVVVVVVVURERFVVVURERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERDMzMzMzMzMzM1VVVVVVVVVVVVVVVURERERERFVVVXd3d3d3d1VVVVVVVXd3d3d3dzMzMzMzM0RERGZmZnd3d2ZmZkRERDMzMyIiIjMzMyIiIiIiIiIiIiIiIhERESIiIiIiIjMzMzMzM0RERFVVVURERDMzMyIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzM0RERDMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERERERERERERERERERDMzM0RERERERFVVVURERERERERERERERFVVVVVVVWZmZmZmZmZmZmZmZmZmZlVVVVVVVURERERERERERERERFVVVWZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZnd3d3d3d2ZmZlVVVURERERERDMzMzMzMzMzM2ZmZmZmZmZmZnd3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiHd3d2ZmZkRERERERERERGZmZmZmZnd3d1VVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVURERERERERERERERFVVVURERERERERERFVVVWZmZlVVVVVVVVVVVWZmZlVVVWZmZkRERERERDMzM0RERDMzM0RERERERERERERERERERFVVVVVVVWZmZlVVVWZmZnd3d4iIiJmZmYiIiGZmZmZmZmZmZlVVVVVVVWZmZlVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERDMzMzMzM0RERERERGZmZmZmZkRERERERDMzM0RERDMzM0RERERERERERERERERERFVVVURERERERDMzM0RERDMzMyIiIkRERERERERERERERERERFVVVURERERERFVVVURERERERDMzM0RERERERFVVVVVVVURERFVVVURERERERDMzMzMzMzMzM1VVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d2ZmZmZmZmZmZnd3d4iIiHd3d2ZmZnd3d4iIiGZmZlVVVVVVVURERERERERERGZmZmZmZlVVVURERFVVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERERERDMzMyIiIjMzM0RERERERERERERERFVVVWZmZmZmZmZmZlVVVVVVVVVVVURERFVVVURERERERDMzM0RERDMzM0RERERERERERDMzMzMzM1VVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVWZmZlVVVVVVVURERERERERERGZmZlVVVVVVVURERERERFVVVVVVVVVVVVVVVURERERERERERERERERERFVVVURERERERFVVVVVVVURERERERERERFVVVVVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVURERERERERERERERFVVVVVVVURERERERDMzMzMzM0RERDMzM0RERDMzMzMzM1VVVWZmZmZmZlVVVWZmZnd3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERERERGZmZmZmZlVVVVVVVVVVVURERERERERERFVVVVVVVVVVVURERFVVVURERERERERERDMzMzMzMyIiIiIiIjMzM1VVVURERERERFVVVVVVVURERERERERERDMzM0RERDMzM0RERERERDMzM0RERDMzM0RERERERERERERERERERERERFVVVWZmZlVVVVVVVURERERERERERERERERERERERERERERERERERERERERERERERERERERERFVVVURERFVVVURERERERERERFVVVURERFVVVURERERERDMzM0RERFVVVVVVVURERERERFVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVURERERERERERERERERERDMzM0RERERERFVVVWZmZmZmZlVVVVVVVURERDMzMzMzMzMzM0RERDMzM0RERERERERERHd3d2ZmZkRERFVVVURERDMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMyIiIjMzMzMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzMyIiIiIiIjMzMzMzMzMzMyIiIjMzMzMzMyIiIiIiIiIiIjMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERERERERERDMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMyIiIiIiIjMzMyIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMyIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzM0RERERERDMzMzMzMzMzMzMzM0RERERERERERDMzMzMzM0RERGZmZlVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVXd3d3d3d5mZmaqqqru7u7u7u7u7u8zMzO7u7v///////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////u7u7d3d3d3d3u7u7d3d3u7u7u7u7u7u7d3d3u7u7d3d3u7u7d3d3u7u7d3d3d3d3u7u7d3d3u7u7u7u7u7u7d3d3u7u7d3d3u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3u7u7MzMzd3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3d3d3MzMzd3d3MzMzMzMzMzMy7u7u7u7u7u7uqqqqqqqqqqqqZmZmqqqqZmZmZmZmZmZmZmZmqqqqqqqqqqqq7u7uqqqq7u7vMzMzMzMzMzMzMzMzd3d3MzMzd3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7u7u7vMzMzMzMzMzMzMzMzMzMzd3d3MzMzd3d3MzMzMzMzMzMy7u7vMzMy7u7uqqqq7u7uqqqq7u7u7u7uqqqq7u7u7u7uqqqqZmZmZmZmZmZmIiIiIiIiIiIh3d3eIiIiIiIiIiIh3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZmZmZmZmZmZmZmIiIiIiIiIiIiIiIh3d3dmZmZmZmZ3d3dmZmZ3d3d3d3eIiIiIiIiIiIiIiIiIiIiZmZmZmZmqqqqZmZmZmZmqqqqqqqqZmZmZmZmZmZmZmZmIiIhmZmZmZmZmZmZVVVVERERERERERERERERERERERERERERERERERERVVVVVVVVERERVVVVVVVVmZmZVVVVERERmZmZ3d3eIiIiqqqq7u7vd3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7u7u7d3d3d3d3u7u7d3d3u7u7u7u7d3d3u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7d3d3d3d3d3d3d3d3u7u7d3d3d3d3u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMzMzMy7u7uqqqqqqqqIiIh3d3d3d3dmZmZVVVVVVVVEREQzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNVVVVmZmZmZmZ3d3dmZmZmZmZmZmZmZmZ3d3d3d3dmZmZ3d3dmZmZVVVVERERERERERERERERVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIREREREREiIiIiIiIiIiIzMzMzMzNERERVVVVVVVVEREQzMzMiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiJEREQzMzNEREREREQiIiIzMzMzMzMzMzNERERERERERERVVVVVVVVVVVVVVVVVVVVERERVVVVERERERERERERVVVVERERVVVVERERERERVVVVERERVVVVmZmZmZmZmZmZmZmZmZmZVVVVEREREREQzMzMzMzNERERmZmZ3d3dmZmZVVVVVVVVmZmZmZmZVVVVmZmZmZmZVVVVmZmZEREREREREREQzMzMiIiIzMzNVVVVmZmZ3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIh3d3dmZmZERERERERVVVVVVVVmZmZ3d3dmZmZmZmZVVVVVVVVERERVVVVVVVVmZmZmZmZVVVVERERERERERERERERERERERERERERERERERERVVVVVVVVVVVVmZmZmZmZmZmZEREREREQzMzMzMzNEREREREREREQzMzMzMzNERERVVVVERERVVVVVVVVVVVVmZmZ3d3d3d3eIiIiZmZl3d3dmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVEREQzMzMzMzNERERERERmZmZVVVVVVVVEREREREREREREREREREREREREREREREREREREREREREREREREREREREQzMzMzMzMzMzNERERERERVVVVERERERERmZmZVVVVERERVVVVERERERERERERVVVVVVVVVVVVEREREREREREREREQzMzMzMzNERERVVVVmZmZERERmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmaIiIiIiIiIiIh3d3dmZmZ3d3dmZmZVVVVVVVVERERERERERERVVVVmZmZVVVVVVVVVVVVVVVVERERERERmZmZVVVVVVVVVVVVVVVVVVVVEREREREREREREREREREREREQzMzMiIiIzMzNERERVVVVERERVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVERERVVVVVVVVEREREREREREREREREREREREQzMzMzMzMzMzNERERVVVVVVVVVVVVmZmZmZmZVVVV3d3dmZmZmZmZmZmZVVVVERERmZmZVVVVVVVVVVVVERERERERERERVVVVERERVVVVERERVVVVERERVVVVmZmZVVVVVVVVERERVVVVERERERERERERERERERERERERVVVVERERVVVVERERERERmZmZVVVVmZmZVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERERERVVVUzMzMzMzMzMzNERERVVVVVVVVEREREREREREREREQzMzNERERVVVUzMzNERERVVVVVVVVmZmZmZmZmZmZ3d3dmZmZ3d3d3d3dmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVVVVVVVVVEREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERmZmZmZmZERERVVVVEREREREREREREREREREREREQzMzNEREQzMzNEREREREQzMzNERERERERERERERERVVVVmZmZmZmZVVVUzMzNEREQzMzNEREQzMzNERERERERERERERERERERERERERERVVVVERERERERVVVVERERERERERERERERERERERERVVVVERERERERERERERERERERVVVVEREREREREREREREREREQzMzMzMzMzMzMzMzMzMzNEREQzMzNERERERERERERERERERERERERERERERERERERERERVVVVmZmZmZmZmZmZVVVVEREQzMzNEREQzMzNEREQzMzNERERERERVVVVERER3d3dmZmZVVVVVVVVEREQzMzMiIiIiIiIzMzMzMzNEREQzMzMzMzNEREREREQzMzMzMzMiIiIzMzMzMzNEREQzMzMzMzNVVVVEREQiIiIiIiIzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzMiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIzMzMiIiIzMzMzMzMzMzMiIiIiIiIzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzNEREREREQzMzMzMzMzMzMzMzNERERVVVVmZmZmZmZmZmZVVVVmZmZVVVVVVVVVVVVmZmZ3d3eIiIiZmZmqqqq7u7vMzMy7u7vMzMzu7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d7u7u3d3d7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMu7u7u7u7qqqqqqqqqqqqmZmZqqqqqqqqmZmZmZmZmZmZmZmZqqqqmZmZqqqqu7u7u7u7zMzMzMzMzMzMzMzM3d3dzMzMzMzM3d3dzMzMzMzMzMzMu7u7zMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7zMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7u7u7qqqqu7u7qqqqu7u7qqqqqqqqmZmZmZmZiIiIiIiIiIiId3d3d3d3d3d3ZmZmd3d3ZmZmd3d3d3d3ZmZmd3d3iIiIiIiIiIiIiIiImZmZmZmZiIiIiIiImZmZmZmZiIiIiIiId3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiImZmZmZmZmZmZmZmZmZmZqqqqqqqqmZmZmZmZmZmZiIiIiIiIZmZmZmZmVVVVVVVVREREREREREREREREREREREREREREREREREREZmZmZmZmVVVVVVVVVVVVREREREREREREZmZmd3d3iIiIiIiImZmZqqqqu7u7zMzM3d3d7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u7u7u3d3d7u7u3d3d7u7u3d3d7u7u3d3d7u7u3d3d3d3d7u7u3d3d7u7u7u7u3d3d7u7u3d3d3d3d3d3d3d3dzMzMu7u7zMzMu7u7u7u7qqqqmZmZiIiIZmZmVVVVREREREREREREMzMzMzMzIiIiMzMzIiIiIiIiIiIiMzMzMzMzMzMzREREMzMzMzMzREREMzMzMzMzREREREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREVVVVZmZmd3d3iIiIiIiImZmZmZmZd3d3ZmZmiIiId3d3iIiIiIiIZmZmVVVVVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiERERIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzIiIiMzMzIiIiERERIiIiERERIiIiIiIiIiIiMzMzIiIiMzMzMzMzIiIiIiIiMzMzMzMzREREMzMzMzMzMzMzREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVREREREREVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVREREVVVVREREMzMzMzMzREREZmZmZmZmVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREMzMzIiIiMzMzZmZmd3d3d3d3d3d3iIiId3d3d3d3iIiImZmZiIiIZmZmd3d3ZmZmd3d3ZmZmVVVVVVVVREREVVVVZmZmiIiId3d3VVVVZmZmVVVVVVVVREREVVVVVVVVREREREREREREREREREREREREVVVVREREREREREREREREVVVVVVVVVVVVVVVVZmZmZmZmVVVVREREMzMzREREREREREREREREREREMzMzREREREREREREVVVVVVVVVVVVZmZmd3d3d3d3d3d3mZmZiIiId3d3ZmZmd3d3ZmZmVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVREREREREREREREREVVVVZmZmVVVVVVVVVVVVVVVVREREREREMzMzREREMzMzREREREREREREMzMzMzMzMzMzREREMzMzMzMzMzMzREREVVVVREREREREVVVVVVVVZmZmREREVVVVVVVVVVVVREREZmZmVVVVVVVVREREMzMzREREMzMzMzMzMzMzMzMzVVVVZmZmVVVVZmZmZmZmVVVVZmZmd3d3d3d3iIiIiIiIiIiIiIiIiIiId3d3ZmZmZmZmZmZmVVVVZmZmVVVVREREREREVVVVZmZmVVVVZmZmVVVVVVVVZmZmVVVVZmZmZmZmd3d3ZmZmVVVVVVVVREREMzMzREREREREMzMzREREREREIiIiMzMzREREVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVREREVVVVREREMzMzREREREREREREREREREREMzMzMzMzMzMzREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmVVVVREREVVVVREREVVVVVVVVREREREREREREREREREREREREVVVVZmZmREREREREREREREREVVVVREREREREREREREREREREREREREREVVVVREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREREREREREVVVVREREREREMzMzIiIiIiIiREREZmZmZmZmVVVVREREREREREREREREREREREREVVVVREREVVVVVVVVZmZmd3d3ZmZmd3d3d3d3ZmZmZmZmZmZmZmZmVVVVREREZmZmVVVVVVVVREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVREREREREVVVVVVVVREREMzMzMzMzREREMzMzMzMzMzMzMzMzREREMzMzREREREREREREZmZmVVVVVVVVVVVVREREREREREREREREREREMzMzREREMzMzREREREREREREREREREREREREVVVVVVVVVVVVVVVVZmZmVVVVREREREREREREREREMzMzREREREREREREREREREREVVVVREREREREREREREREVVVVREREREREREREREREREREREREREREREREREREREREMzMzREREZmZmZmZmVVVVREREREREREREMzMzMzMzREREREREREREREREREREMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzREREVVVVVVVVVVVVZmZmVVVVREREREREMzMzMzMzREREREREREREREREREREREREZmZmiIiIZmZmVVVVVVVVREREMzMzMzMzMzMzIiIiMzMzREREIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREVVVVMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiIiIiMzMzIiIiMzMzIiIiIiIiMzMzIiIiMzMzMzMzREREREREMzMzREREREREREREREREIiIiMzMzMzMzMzMzMzMzIiIiMzMzREREREREIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREVVVVVVVVd3d3d3d3ZmZmVVVVVVVVZmZmd3d3d3d3iIiImZmZqqqqu7u7zMzMzMzMzMzM7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////+7u7v///////+7u7v///+7u7v///+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3d3d3e7u7t3d3d3d3czMzN3d3czMzN3d3d3d3e7u7t3d3d3d3d3d3czMzN3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzLu7u7u7u6qqqqqqqqqqqqqqqpmZmaqqqpmZmaqqqqqqqqqqqqqqqqqqqru7u7u7u7u7u7u7u7u7u8zMzLu7u8zMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u8zMzLu7u8zMzLu7u8zMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u6qqqqqqqpmZmZmZmYiIiIiIiHd3d3d3d3d3d2ZmZlVVVWZmZmZmZlVVVWZmZlVVVWZmZnd3d2ZmZnd3d4iIiJmZmYiIiIiIiIiIiJmZmZmZmZmZmZmZmYiIiIiIiIiIiHd3d3d3d2ZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d4iIiHd3d4iIiIiIiJmZmZmZmZmZmaqqqqqqqpmZmYiIiIiIiJmZmXd3d2ZmZlVVVWZmZmZmZkRERERERERERERERERERERERGZmZlVVVVVVVVVVVVVVVURERERERDMzMzMzMzMzMzMzM0RERFVVVWZmZoiIiKqqqszMzN3d3d3d3d3d3d3d3d3d3e7u7u7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7v///+7u7u7u7u7u7v///+7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3e7u7t3d3d3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7u7u7t3d3e7u7t3d3d3d3d3d3d3d3czMzLu7u7u7u6qqqpmZmZmZmXd3d3d3d2ZmZmZmZmZmZlVVVVVVVURERERERERERERERERERERERERERDMzM0RERFVVVVVVVWZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVURERERERERERERERDMzMzMzM0RERFVVVVVVVVVVVXd3d4iIiIiIiIiIiKqqqoiIiHd3d3d3d5mZmYiIiJmZmZmZmWZmZlVVVURERDMzMzMzM0RERDMzMzMzMyIiIiIiIiIiIiIiIhERESIiIiIiIiIiIhERESIiIiIiIhERESIiIhERERERESIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIjMzMyIiIjMzMyIiIjMzM0RERERERDMzM0RERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERDMzM0RERERERFVVVVVVVURERERERFVVVVVVVVVVVVVVVWZmZlVVVVVVVURERERERERERDMzM0RERDMzM0RERERERFVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVURERFVVVTMzM0RERERERGZmZnd3d3d3d2ZmZnd3d2ZmZmZmZnd3d3d3d3d3d3d3d2ZmZkRERFVVVVVVVVVVVURERFVVVVVVVWZmZnd3d4iIiHd3d2ZmZmZmZlVVVWZmZmZmZlVVVURERERERERERFVVVVVVVURERERERDMzM0RERERERERERERERFVVVVVVVWZmZmZmZmZmZmZmZlVVVURERERERERERFVVVTMzM0RERDMzM0RERERERERERERERERERFVVVVVVVWZmZnd3d4iIiIiIiHd3d2ZmZnd3d2ZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVURERDMzM0RERERERFVVVWZmZlVVVVVVVVVVVVVVVURERERERERERDMzM0RERDMzM0RERERERERERDMzMzMzMzMzMzMzMzMzM0RERGZmZmZmZlVVVURERGZmZmZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVTMzM0RERDMzMzMzMzMzMzMzMzMzM1VVVWZmZmZmZmZmZnd3d2ZmZmZmZnd3d3d3d3d3d3d3d4iIiIiIiHd3d2ZmZmZmZmZmZlVVVVVVVVVVVWZmZkRERERERFVVVXd3d2ZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZnd3d3d3d1VVVURERERERERERERERERERERERERERDMzMzMzMzMzM0RERGZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVURERERERERERDMzMzMzM0RERERERDMzM1VVVTMzMzMzM0RERDMzM0RERFVVVVVVVWZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZnd3d1VVVURERFVVVVVVVURERERERERERERERERERFVVVURERERERERERFVVVURERERERERERERERERERERERFVVVURERERERERERERERERERERERFVVVURERFVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzM1VVVWZmZmZmZkRERERERDMzMzMzM0RERERERERERERERERERGZmZnd3d4iIiHd3d2ZmZnd3d3d3d2ZmZlVVVVVVVURERFVVVVVVVURERERERERERFVVVURERFVVVURERFVVVURERFVVVVVVVVVVVWZmZlVVVURERFVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERDMzM0RERERERFVVVVVVVVVVVURERFVVVVVVVURERERERERERERERDMzM0RERERERERERERERERERERERFVVVVVVVURERERERFVVVWZmZmZmZlVVVURERERERERERERERERERERERERERERERERERERERFVVVWZmZmZmZlVVVURERFVVVURERERERERERERERERERERERERERERERERERFVVVURERGZmZnd3d2ZmZlVVVURERERERERERDMzMzMzM0RERERERERERERERDMzM0RERERERDMzM0RERDMzM0RERERERFVVVVVVVURERFVVVVVVVVVVVURERERERERERERERERERERERFVVVURERERERFVVVWZmZmZmZlVVVVVVVURERFVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM0RERERERDMzMzMzMyIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERDMzM0RERERERERERERERDMzMyIiIjMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIjMzM0RERDMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIhERESIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMyIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERERERGZmZnd3d3d3d2ZmZlVVVWZmZnd3d3d3d4iIiIiIiJmZmaqqqru7u7u7u8zMzO7u7v///+7u7v///////////////////+7u7v///////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////u7u7u7u7////u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3u7u7d3d3d3d3u7u7u7u7u7u7d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7uqqqqqqqqqqqqqqqqqqqqZmZmqqqqqqqqZmZmqqqqZmZmqqqqqqqqqqqqqqqq7u7u7u7u7u7u7u7u7u7vMzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7uqqqq7u7u7u7u7u7u7u7u7u7u7u7vMzMy7u7u7u7u7u7u7u7uqqqq7u7uqqqqqqqqZmZmZmZmZmZmIiIh3d3eIiIh3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZVVVVmZmZmZmZmZmZ3d3eIiIiIiIiIiIiZmZmqqqqZmZmZmZmZmZmZmZmZmZmIiIh3d3dmZmZVVVV3d3d3d3d3d3d3d3dmZmZ3d3dmZmZmZmZmZmZ3d3d3d3d3d3d3d3eZmZmqqqqZmZmqqqqqqqqZmZmIiIh3d3d3d3d3d3dVVVVVVVVVVVVERERERERERERERERmZmZVVVVVVVVmZmZVVVVVVVVVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzNVVVVmZmaIiIiZmZmqqqrMzMzd3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7////u7u7u7u7////u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3u7u7d3d3d3d3d3d3d3d3u7u7d3d3u7u7d3d3u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3MzMy7u7u7u7uqqqqqqqqZmZmZmZmIiIiIiIiIiIh3d3d3d3d3d3d3d3dmZmZ3d3d3d3dmZmZ3d3dmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmaIiIiIiIiIiIh3d3d3d3d3d3d3d3dmZmZmZmZmZmZVVVVVVVVVVVVEREQzMzNERERERERERERVVVVVVVVmZmZ3d3d3d3d3d3eIiIiqqqqZmZl3d3eZmZmZmZmIiIiIiIh3d3d3d3dmZmZEREQzMzNEREQzMzMzMzMiIiIiIiIREREiIiIiIiIREREREREREREREREiIiIiIiIiIiIiIiIREREiIiIiIiIREREiIiIzMzMiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNERERERERVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVEREREREQzMzMzMzNERERVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZVVVVVVVVEREREREQzMzNEREQzMzNERERERERVVVV3d3dmZmZVVVVVVVVVVVVERERVVVVmZmZVVVVmZmZVVVVVVVVERERERERERERERERVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVmZmZ3d3d3d3dmZmZVVVVVVVVVVVVEREREREQzMzNERERVVVVVVVVmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVERERERERVVVVVVVVVVVVERERERERERERERERVVVVVVVVERERVVVVmZmZ3d3dmZmZmZmZVVVVERERERERVVVUzMzNERERERERERERERERERERERERERERVVVVVVVVmZmZmZmZmZmaIiIiIiIhmZmZVVVVmZmZmZmZmZmZ3d3dmZmZVVVVVVVVmZmZmZmZVVVVmZmZmZmZmZmZVVVVmZmZmZmZVVVVVVVVERERERERERERVVVVmZmZVVVVVVVVERERERERVVVVEREQzMzNERERERERERERmZmZmZmZVVVVEREQzMzMzMzMzMzMzMzNERERVVVVVVVVVVVVVVVVmZmZ3d3dVVVVVVVVVVVVmZmZmZmZmZmZVVVVEREQzMzNEREQzMzMzMzMzMzMzMzMzMzNVVVVVVVVmZmZ3d3dmZmZmZmZmZmZ3d3eIiIiIiIh3d3eIiIiIiIh3d3dmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVERERVVVVmZmZ3d3dVVVVVVVV3d3d3d3dmZmZVVVVmZmaIiIh3d3dEREREREREREQzMzNEREQzMzNEREREREQzMzMzMzMzMzMzMzNVVVV3d3dmZmZVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVEREQzMzNEREQzMzMzMzNEREREREREREREREQzMzNERERERERERERVVVVVVVVVVVVmZmZmZmZVVVVVVVVmZmZmZmZ3d3dmZmZVVVVERERVVVVVVVVEREREREREREQzMzNERERVVVVEREREREREREREREREREQzMzNERERERERERERVVVVERERERERERERVVVUzMzNERERERERVVVVERERVVVVERERERERVVVVERERVVVVEREREREREREREREREREREREREREREREREREREREREREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzNERERVVVVVVVVEREQzMzMzMzMzMzNERERERERERERVVVVmZmZ3d3d3d3d3d3d3d3eIiIh3d3dVVVVERERERERVVVVERERVVVVERERERERERERERERERERVVVVERERERERERERVVVVmZmZ3d3dmZmZVVVVVVVVVVVVEREREREQzMzNEREQzMzMzMzMzMzNEREREREREREREREQzMzNEREQzMzNEREQzMzNERERVVVVERERVVVVVVVVERERVVVVERERERERERERERERERERVVVVERERERERERERERERERERERERVVVVERERmZmZ3d3dVVVVERERVVVVEREREREQzMzNEREQzMzNERERVVVVmZmZVVVVmZmZmZmZERERVVVVVVVVEREREREQzMzNERERERERERERERERERERERERERERVVVV3d3eIiIhmZmZmZmZEREREREREREREREREREREREREREQzMzNEREREREQzMzNEREREREQzMzNERERVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERVVVVERERERERVVVVVVVVVVVVEREREREQzMzNEREREREREREQzMzNEREREREQzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzMzMzNEREREREQzMzMiIiIzMzMiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzNEREQzMzNERERERERVVVVEREQzMzMzMzMiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzNEREQzMzMzMzMzMzMzMzMiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIzMzMzMzMiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVmZmZ3d3dmZmZVVVVmZmZ3d3d3d3d3d3eIiIiIiIiZmZmZmZm7u7u7u7u7u7vd3d3///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u7u7u3d3d7u7u3d3d7u7u3d3d7u7u3d3d7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3dzMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3dzMzM3d3d3d3dzMzMzMzMzMzMu7u7u7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqqqqqmZmZmZmZmZmZmZmZqqqqqqqqmZmZqqqqu7u7u7u7zMzMzMzMu7u7zMzM3d3dzMzMzMzMu7u7u7u7u7u7qqqqqqqqu7u7qqqqqqqqqqqqqqqqqqqqu7u7u7u7u7u7qqqqu7u7qqqqu7u7qqqqqqqqqqqqmZmZmZmZmZmZiIiIiIiId3d3ZmZmZmZmd3d3ZmZmd3d3d3d3d3d3d3d3ZmZmZmZmVVVVZmZmZmZmZmZmd3d3iIiImZmZmZmZmZmZqqqqqqqqqqqqmZmZmZmZmZmZmZmZiIiId3d3d3d3iIiIZmZmd3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmVVVVd3d3iIiIiIiImZmZmZmZmZmZmZmZmZmZiIiIiIiIZmZmZmZmVVVVZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVMzMzMzMzMzMzMzMzMzMzREREREREVVVVVVVVd3d3mZmZu7u7zMzM7u7u////7u7u7u7u7u7u7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d3d3d7u7u3d3dzMzMzMzMzMzMu7u7qqqqqqqqqqqqmZmZmZmZmZmZmZmZiIiImZmZmZmZmZmZiIiId3d3d3d3iIiId3d3iIiIiIiId3d3mZmZmZmZmZmZiIiIiIiId3d3d3d3d3d3iIiId3d3d3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVREREREREREREREREMzMzREREREREVVVVVVVVVVVVZmZmd3d3iIiIiIiId3d3iIiIqqqqd3d3ZmZmZmZmd3d3ZmZmREREREREMzMzREREMzMzIiIiIiIiERERIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVVVVVZmZmZmZmZmZmVVVVZmZmd3d3ZmZmVVVVREREREREMzMzMzMzMzMzVVVVVVVVZmZmVVVVVVVVVVVVZmZmZmZmd3d3ZmZmREREMzMzMzMzREREVVVVVVVVREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmVVVVVVVVREREREREMzMzREREREREVVVVREREREREZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmVVVVVVVVREREVVVVVVVVREREREREREREVVVVVVVVZmZmd3d3d3d3ZmZmd3d3ZmZmVVVVREREVVVVREREREREREREVVVVVVVVREREVVVVVVVVREREVVVVREREREREVVVVd3d3iIiIZmZmREREVVVVREREREREMzMzREREVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVVVVVZmZmd3d3qqqqiIiIZmZmZmZmd3d3ZmZmZmZmZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmREREVVVVVVVVZmZmZmZmZmZmVVVVREREREREREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVREREREREMzMzMzMzREREVVVVREREVVVVVVVVVVVVZmZmd3d3ZmZmVVVVZmZmZmZmd3d3ZmZmREREREREMzMzREREREREMzMzMzMzMzMzMzMzREREVVVVZmZmZmZmd3d3d3d3d3d3d3d3iIiIiIiIiIiId3d3iIiId3d3VVVVZmZmVVVVZmZmREREREREREREVVVVREREREREVVVVZmZmVVVVZmZmd3d3d3d3ZmZmVVVVZmZmd3d3ZmZmVVVVREREREREMzMzREREMzMzREREMzMzMzMzMzMzMzMzMzMzREREZmZmZmZmVVVVVVVVZmZmVVVVVVVVVVVVREREREREREREMzMzREREMzMzREREREREREREREREREREREREREREREREREREREREZmZmZmZmZmZmZmZmVVVVZmZmZmZmVVVVVVVVVVVVREREREREVVVVVVVVREREREREREREREREREREREREREREMzMzREREREREREREREREREREREREREREVVVVREREREREVVVVVVVVMzMzREREREREVVVVREREREREVVVVVVVVREREVVVVREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREMzMzMzMzREREMzMzMzMzMzMzREREREREREREREREMzMzMzMzMzMzREREREREREREVVVVZmZmZmZmd3d3iIiIiIiIiIiIZmZmVVVVREREREREVVVVREREVVVVREREVVVVREREREREREREREREREREREREREREVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREMzMzMzMzREREREREREREREREREREREREREREMzMzREREREREMzMzREREREREREREVVVVVVVVVVVVVVVVREREREREREREREREREREVVVVVVVVREREREREREREREREREREREREVVVVREREVVVVZmZmZmZmVVVVVVVVVVVVREREREREMzMzREREREREVVVVZmZmVVVVREREREREZmZmVVVVVVVVVVVVREREREREREREREREREREREREREREREREVVVVVVVVd3d3iIiIZmZmZmZmZmZmREREMzMzREREREREREREREREREREREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREVVVVVVVVVVVVVVVVREREVVVVREREREREVVVVREREVVVVVVVVREREREREMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREREREMzMzMzMzREREREREMzMzREREMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzREREREREVVVVREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzREREMzMzREREREREMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzIiIiIiIiMzMzREREMzMzMzMzREREVVVVVVVVZmZmd3d3ZmZmd3d3d3d3VVVVd3d3iIiIiIiIiIiIqqqqqqqqqqqqzMzM7u7u7u7u////7u7u////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3e7u7t3d3e7u7t3d3e7u7u7u7u7u7t3d3e7u7u7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7t3d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzLu7u8zMzLu7u8zMzMzMzMzMzMzMzMzMzN3d3czMzMzMzMzMzN3d3czMzN3d3czMzN3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u6qqqqqqqqqqqqqqqqqqqpmZmaqqqqqqqqqqqqqqqru7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqru7u6qqqqqqqqqqqpmZmaqqqpmZmZmZmaqqqpmZmaqqqpmZmaqqqqqqqqqqqqqqqru7u6qqqqqqqqqqqqqqqpmZmYiIiHd3d3d3d3d3d2ZmZmZmZmZmZlVVVWZmZnd3d3d3d2ZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZmZmZnd3d5mZmYiIiJmZmZmZmZmZmaqqqqqqqoiIiHd3d4iIiIiIiHd3d3d3d3d3d2ZmZlVVVVVVVVVVVTMzM1VVVWZmZmZmZmZmZmZmZoiIiIiIiIiIiJmZmZmZmYiIiHd3d3d3d4iIiGZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZlVVVURERDMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzM1VVVWZmZpmZmaqqqru7u8zMzN3d3d3d3d3d3e7u7t3d3e7u7u7u7t3d3e7u7t3d3e7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7t3d3e7u7u7u7u7u7t3d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3czMzLu7u7u7u6qqqpmZmZmZmZmZmZmZmZmZmZmZmaqqqqqqqpmZmYiIiJmZmYiIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiJmZmZmZmZmZmZmZmZmZmZmZmYiIiHd3d3d3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d2ZmZlVVVVVVVVVVVURERERERERERERERERERFVVVURERFVVVWZmZoiIiIiIiIiIiGZmZlVVVYiIiJmZmXd3d2ZmZmZmZlVVVVVVVURERERERERERDMzMyIiIiIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERDMzM1VVVWZmZnd3d3d3d2ZmZnd3d3d3d3d3d2ZmZmZmZlVVVURERDMzMzMzM1VVVVVVVWZmZlVVVURERFVVVVVVVWZmZnd3d2ZmZlVVVURERERERFVVVVVVVVVVVVVVVURERERERERERGZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZkRERDMzMzMzM0RERERERERERDMzM1VVVVVVVWZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d3d3d1VVVVVVVVVVVURERERERFVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVURERDMzM1VVVWZmZmZmZlVVVVVVVVVVVURERDMzM0RERERERFVVVURERERERERERFVVVWZmZlVVVVVVVVVVVWZmZoiIiJmZmYiIiIiIiGZmZnd3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVWZmZnd3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZkRERERERERERERERCIiIjMzM1VVVWZmZlVVVVVVVWZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVURERERERERERDMzMzMzMzMzMzMzMzMzM0RERERERGZmZmZmZmZmZmZmZnd3d3d3d3d3d2ZmZnd3d3d3d3d3d2ZmZmZmZlVVVVVVVVVVVURERERERERERFVVVVVVVURERFVVVWZmZlVVVWZmZmZmZnd3d3d3d1VVVVVVVVVVVVVVVURERERERERERERERERERDMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM1VVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVURERFVVVURERDMzMzMzMzMzM0RERERERFVVVVVVVURERERERERERERERDMzM0RERGZmZnd3d2ZmZmZmZlVVVVVVVVVVVURERERERERERERERERERERERERERFVVVVVVVURERDMzMzMzMzMzM1VVVURERDMzMzMzM0RERERERDMzM0RERERERERERERERFVVVVVVVURERERERERERERERERERFVVVURERFVVVURERERERERERERERERERERERERERERERERERERERFVVVURERERERERERFVVVURERDMzM0RERDMzM0RERERERDMzM0RERERERERERERERERERDMzMzMzMzMzM0RERDMzMzMzM0RERERERFVVVVVVVXd3d3d3d3d3d2ZmZlVVVURERERERERERFVVVVVVVVVVVURERERERERERERERERERERERERERERERERERFVVVURERFVVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERDMzM0RERERERERERERERERERERERDMzM0RERERERFVVVVVVVVVVVURERERERFVVVURERFVVVURERFVVVURERERERERERERERERERFVVVURERERERFVVVVVVVWZmZlVVVVVVVVVVVURERERERERERERERERERERERFVVVTMzM0RERFVVVVVVVVVVVVVVVURERERERERERERERERERERERFVVVURERFVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVURERERERERERFVVVVVVVURERFVVVURERERERERERFVVVYiIiIiIiGZmZlVVVURERERERERERERERERERERERERERERERERERFVVVURERERERFVVVURERERERERERERERERERCIiIjMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERERERERERDMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzMyIiIjMzMyIiIjMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVURERERERDMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzM0RERERERDMzMzMzM0RERERERERERERERERERERERDMzM0RERDMzMzMzM0RERDMzMzMzM0RERERERERERDMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMzMzM0RERERERDMzMzMzM0RERDMzMzMzM0RERDMzMzMzMzMzMyIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVWZmZmZmZnd3d2ZmZmZmZnd3d4iIiJmZmZmZmZmZmaqqqpmZmaqqqru7u93d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////u7u7u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3u7u7d3d3d3d3u7u7d3d3u7u7d3d3u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMy7u7u7u7vMzMzMzMzMzMy7u7u7u7u7u7vMzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMy7u7vMzMzMzMzMzMy7u7uqqqqqqqqqqqqqqqqqqqqqqqqqqqq7u7u7u7uqqqq7u7uqqqq7u7uqqqqqqqqqqqqqqqqqqqqqqqqqqqqZmZmqqqqZmZmqqqqZmZmqqqqZmZmqqqqqqqqZmZmZmZmZmZmZmZmqqqqZmZmqqqqqqqqqqqqqqqq7u7uqqqqZmZmZmZmZmZmIiIh3d3dmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3eIiIiZmZmZmZmZmZmIiIiIiIiZmZmZmZmZmZmIiIiIiIh3d3dmZmZmZmZERERVVVVVVVV3d3dmZmZERERVVVV3d3d3d3dmZmZmZmZ3d3dmZmaIiIiIiIiIiIh3d3d3d3d3d3d3d3dmZmZ3d3d3d3dmZmZmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVVEREREREREREQzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNERERERERVVVVmZmZ3d3eZmZmqqqq7u7vd3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3MzMy7u7uqqqq7u7uZmZmqqqqqqqqIiIiIiIiIiIiZmZmIiIiIiIiIiIiZmZmIiIiIiIh3d3d3d3d3d3d3d3dmZmZmZmZVVVVERERmZmZ3d3eIiIiIiIiZmZmIiIh3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3eIiIh3d3d3d3dmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3eIiIiIiIiZmZmqqqrMzMzu7u7d3d27u7tmZmZVVVVVVVV3d3d3d3dmZmZmZmZEREREREREREREREQzMzMiIiIiIiIiIiIREREREREiIiIiIiIiIiIiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIREREiIiIiIiIzMzMzMzMzMzMiIiIiIiIzMzMiIiIzMzMzMzNEREREREQzMzMzMzNVVVVERERERERERERERERVVVVmZmZmZmZ3d3d3d3dmZmZmZmZmZmZmZmZmZmZEREQzMzMzMzNVVVVmZmZmZmZVVVVERERERERERERVVVVmZmZ3d3dVVVVERERVVVVERERERERERERERERERERERERERERVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVEREREREREREQzMzNERERERERERERERERVVVVmZmZmZmZmZmZ3d3d3d3dmZmZmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVERERVVVV3d3d3d3d3d3dmZmZVVVVVVVVVVVVERERERERERERVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVEREREREQzMzNERERVVVVmZmZmZmZVVVVERERERERERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZ3d3eZmZl3d3eIiIh3d3d3d3eIiIhmZmZmZmZmZmZ3d3dmZmZmZmZ3d3eIiIiIiIiIiIiZmZl3d3d3d3dmZmZmZmZVVVVVVVVmZmZ3d3dmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVEREREREREREQzMzMiIiIzMzNERERmZmZmZmZVVVVmZmZmZmZmZmZ3d3dmZmZVVVVmZmZVVVVEREREREQzMzNEREREREQzMzMzMzMzMzNERERERERVVVVERERmZmZ3d3dmZmZmZmZ3d3d3d3d3d3dmZmZ3d3dmZmZmZmZmZmZmZmZERERVVVVVVVVERERERERVVVVVVVVVVVVERERERERmZmZ3d3dVVVVVVVVVVVVmZmZVVVVVVVVVVVVERERERERERERERERERERERERVVVVEREREREQzMzMzMzMzMzMzMzMiIiJERER3d3dmZmZVVVVmZmZmZmZVVVVERERERERVVVVEREREREREREQzMzNVVVVVVVVmZmZVVVVEREREREQzMzMzMzMzMzNERERVVVVVVVVmZmZmZmZVVVVEREREREQzMzNEREREREQzMzNERERERERVVVVVVVVVVVVEREREREQzMzMzMzNEREREREREREREREQzMzMzMzNERERERERERERVVVVmZmZVVVVEREREREREREREREQzMzNERERERERVVVVERERERERVVVVERERERERVVVVERERERERERERERERERERVVVVEREREREREREREREQzMzNEREQzMzNEREREREREREQzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNERERERERmZmZ3d3d3d3dVVVVVVVVERERVVVVERERVVVVVVVVVVVVEREREREREREREREREREREREREREQzMzNERERERERERERERERERERVVVVVVVVVVVVERERERERERERVVVVVVVVVVVVEREREREREREREREREREQzMzNERERERERERERERERERERERERERERVVVVERERERERERERVVVVERERVVVVVVVVVVVVERERERERERERERERERERERERERERERERERERERERERERmZmZVVVVVVVVVVVVEREREREQzMzNEREREREQzMzNERERERERERERERERVVVVmZmZVVVVVVVVERERERERERERERERERERERERVVVVVVVVmZmZVVVVVVVVEREREREQzMzNERERERERVVVVmZmZERERVVVVVVVVVVVVEREREREQzMzNERERmZmZ3d3dEREREREREREREREQzMzNERERERERERERERERERERVVVVVVVVERERVVVVERERVVVVEREREREQzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVEREQzMzNEREQzMzNEREQzMzNEREQzMzMzMzNEREREREQzMzMzMzMzMzMiIiIiIiIzMzNEREQzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNEREQzMzNEREQzMzMzMzNERERERERERERVVVVEREREREQzMzMzMzMzMzMzMzMzMzNERERVVVVEREREREQzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERmZmZmZmZ3d3dmZmaIiIiZmZmZmZmZmZmZmZmZmZmZmZmZmZmqqqrMzMzu7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3dzMzM3d3dzMzMzMzM3d3dzMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzM3d3dzMzMzMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7zMzMu7u7u7u7u7u7zMzMzMzMu7u7zMzMzMzMzMzMzMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzMzMzMu7u7u7u7u7u7u7u7qqqqqqqqqqqqqqqqu7u7qqqqu7u7qqqqu7u7qqqqqqqqqqqqmZmZiIiIiIiIiIiIiIiImZmZmZmZmZmZmZmZmZmZqqqqmZmZqqqqmZmZqqqqmZmZqqqqmZmZmZmZmZmZmZmZmZmZmZmZmZmZqqqqmZmZmZmZqqqqmZmZmZmZmZmZd3d3d3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmd3d3d3d3d3d3d3d3iIiIiIiImZmZiIiImZmZmZmZiIiId3d3ZmZmZmZmVVVVd3d3d3d3ZmZmVVVVVVVVZmZmVVVVREREVVVVVVVVd3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiId3d3ZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREMzMzREREMzMzMzMzMzMzMzMzREREREREVVVVREREREREREREREREVVVViIiImZmZu7u73d3d7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3dzMzMzMzMu7u7qqqqqqqqiIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmVVVVZmZmVVVVVVVVREREREREREREREREVVVVZmZmd3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3iIiId3d3d3d3d3d3ZmZmZmZmVVVVZmZmZmZmd3d3d3d3iIiIqqqqu7u7u7u7zMzM3d3d7u7u7u7u////7u7u7u7uqqqqZmZmREREREREZmZmZmZmZmZmVVVVVVVVMzMzMzMzREREMzMzMzMzIiIiERERIiIiERERIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiIiIiMzMzMzMzIiIiMzMzIiIiIiIiIiIiMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiMzMzREREMzMzREREREREVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmd3d3ZmZmVVVVVVVVREREVVVVREREMzMzREREREREVVVVZmZmd3d3ZmZmREREMzMzREREVVVVVVVVVVVVVVVVREREMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREREREREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVZmZmd3d3ZmZmZmZmZmZmVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREZmZmmZmZd3d3ZmZmVVVVVVVVREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVREREVVVVREREREREZmZmZmZmVVVVREREREREREREREREVVVVREREREREVVVVREREVVVVREREVVVVVVVVZmZmd3d3iIiId3d3d3d3d3d3iIiIiIiId3d3ZmZmZmZmZmZmd3d3d3d3d3d3mZmZiIiImZmZiIiId3d3d3d3ZmZmZmZmREREVVVVZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVREREREREREREREREMzMzIiIiMzMzMzMzZmZmZmZmVVVVVVVVZmZmZmZmd3d3ZmZmZmZmVVVVREREREREMzMzREREREREMzMzMzMzREREREREREREREREREREVVVVVVVVd3d3d3d3ZmZmd3d3d3d3iIiId3d3d3d3VVVVZmZmZmZmVVVVVVVVVVVVREREVVVVREREREREVVVVVVVVVVVVREREVVVVd3d3ZmZmREREVVVVVVVVVVVVREREVVVVREREMzMzREREMzMzVVVVREREVVVVMzMzMzMzMzMzMzMzREREREREMzMzREREVVVVZmZmZmZmZmZmZmZmVVVVREREREREREREREREMzMzREREREREVVVVVVVVZmZmREREVVVVREREMzMzMzMzMzMzREREREREVVVVVVVVVVVVVVVVREREMzMzREREREREMzMzREREVVVVREREVVVVREREREREMzMzMzMzMzMzMzMzREREREREMzMzREREREREREREREREREREVVVVZmZmd3d3VVVVREREMzMzREREREREMzMzREREREREVVVVREREVVVVREREREREREREREREVVVVREREVVVVREREVVVVREREREREMzMzREREREREREREMzMzREREREREREREREREMzMzREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREVVVVZmZmZmZmVVVVVVVVREREREREVVVVVVVVVVVVREREVVVVREREREREREREREREREREREREREREREREREREREREREREREREVVVVZmZmVVVVREREREREREREVVVVREREVVVVREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREVVVVVVVVREREREREVVVVREREZmZmVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREREREREREREREREREVVVVZmZmVVVVREREREREREREVVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVREREMzMzREREVVVVREREVVVVVVVVVVVVVVVVVVVVREREREREMzMzREREMzMzREREMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREREREREREREREREREVVVVREREVVVVMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVVVVVREREMzMzREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzREREREREMzMzIiIiMzMzMzMzMzMzMzMzVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzVVVVZmZmREREMzMzREREMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREREREREREREREMzMzMzMzREREREREREREREREREREREREREREMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzIiIiREREREREREREMzMzMzMzMzMzMzMzREREREREMzMzMzMzMzMzREREMzMzREREMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzREREREREVVVVVVVVZmZmZmZmZmZmd3d3mZmZmZmZmZmZmZmZiIiIiIiIqqqqqqqqqqqqzMzM3d3d7u7u////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////+7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzLu7u7u7u7u7u7u7u6qqqru7u6qqqqqqqqqqqru7u6qqqru7u6qqqru7u7u7u7u7u8zMzMzMzN3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3czMzN3d3czMzN3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u8zMzLu7u7u7u8zMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u8zMzMzMzMzMzN3d3czMzN3d3czMzN3d3czMzMzMzMzMzLu7u6qqqru7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqpmZmXd3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiJmZmaqqqoiIiJmZmZmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiJmZmYiIiIiIiIiIiKqqqpmZmZmZmZmZmYiIiIiIiIiIiHd3d2ZmZmZmZmZmZlVVVURERERERERERERERFVVVURERFVVVURERGZmZlVVVVVVVVVVVVVVVVVVVWZmZnd3d2ZmZoiIiIiIiJmZmYiIiIiIiIiIiIiIiIiIiHd3d4iIiIiIiHd3d2ZmZlVVVVVVVURERERERFVVVVVVVWZmZlVVVWZmZnd3d3d3d2ZmZmZmZnd3d4iIiIiIiIiIiHd3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVURERDMzMzMzM0RERERERERERFVVVURERERERERERDMzM0RERFVVVWZmZpmZmbu7u8zMzN3d3d3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3czMzKqqqpmZmYiIiIiIiHd3d3d3d2ZmZnd3d3d3d3d3d4iIiHd3d3d3d3d3d3d3d2ZmZmZmZkRERERERFVVVWZmZnd3d4iIiJmZmaqqqpmZmaqqqpmZmYiIiHd3d2ZmZnd3d3d3d2ZmZmZmZnd3d4iIiJmZmaqqqru7u8zMzN3d3d3d3e7u7u7u7u7u7v///+7u7t3d3czMzMzMzKqqqoiIiGZmZkRERERERERERFVVVVVVVVVVVVVVVURERERERDMzMzMzM0RERDMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzM1VVVVVVVVVVVVVVVWZmZmZmZlVVVWZmZnd3d2ZmZlVVVTMzM0RERERERERERDMzMzMzMzMzM1VVVVVVVWZmZmZmZlVVVURERERERFVVVURERERERERERDMzMzMzMzMzM0RERERERERERDMzM0RERERERFVVVVVVVWZmZmZmZmZmZkRERERERFVVVVVVVVVVVTMzM0RERERERDMzMzMzM0RERERERFVVVVVVVURERERERFVVVWZmZnd3d3d3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVVVVVURERFVVVXd3d3d3d2ZmZmZmZmZmZlVVVURERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVWZmZlVVVVVVVURERERERERERERERERERERERERERERERERERFVVVVVVVWZmZmZmZoiIiHd3d2ZmZnd3d4iIiIiIiHd3d3d3d3d3d3d3d3d3d4iIiIiIiJmZmYiIiJmZmZmZmYiIiIiIiGZmZlVVVVVVVURERFVVVWZmZmZmZoiIiIiIiHd3d4iIiHd3d4iIiGZmZmZmZlVVVWZmZlVVVURERERERERERERERERERDMzMzMzMyIiIjMzM1VVVWZmZlVVVVVVVVVVVXd3d2ZmZmZmZmZmZlVVVURERDMzMzMzMzMzM0RERERERERERERERERERFVVVURERFVVVURERFVVVWZmZnd3d3d3d3d3d2ZmZnd3d3d3d2ZmZmZmZmZmZmZmZlVVVVVVVURERERERFVVVURERERERERERFVVVVVVVURERERERERERGZmZmZmZlVVVVVVVURERERERERERERERDMzMzMzM0RERERERFVVVURERERERDMzMzMzMzMzMzMzM0RERERERERERDMzM0RERFVVVVVVVVVVVURERERERDMzM0RERERERERERERERFVVVURERFVVVVVVVURERERERDMzMzMzMzMzMzMzMzMzM0RERERERFVVVURERFVVVURERDMzMzMzMzMzM0RERERERERERFVVVURERERERERERDMzM0RERERERDMzMzMzMzMzMzMzM0RERFVVVVVVVURERERERFVVVVVVVWZmZlVVVURERDMzM0RERFVVVURERERERERERERERERERERERERERERERERERERERFVVVURERERERERERERERERERERERERERDMzM0RERERERDMzM0RERDMzM0RERERERDMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERGZmZmZmZlVVVVVVVURERERERFVVVVVVVVVVVVVVVURERERERFVVVURERERERERERERERERERERERERERERERERERFVVVVVVVVVVVURERERERERERERERERERFVVVURERDMzMzMzM0RERDMzM0RERERERERERERERERERERERERERERERERERERERERERFVVVWZmZmZmZlVVVVVVVVVVVVVVVURERERERERERFVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERERERDMzMzMzM0RERGZmZmZmZlVVVURERERERFVVVURERFVVVVVVVVVVVWZmZmZmZmZmZkRERERERERERERERERERFVVVURERERERFVVVVVVVURERDMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERERERDMzM0RERERERERERERERERERERERERERERERERERDMzMzMzMzMzMyIiIjMzMyIiIjMzM0RERERERDMzMzMzMzMzM0RERDMzMzMzM1VVVVVVVVVVVURERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMyIiIjMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERFVVVURERDMzMzMzMzMzMzMzMzMzM0RERFVVVURERERERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVURERERERDMzM0RERERERERERERERERERERERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzM0RERFVVVURERDMzMzMzM0RERFVVVVVVVTMzM0RERDMzMzMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIhERERERERERERERESIiIhERESIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIjMzMyIiIjMzMzMzM0RERERERFVVVVVVVWZmZnd3d2ZmZmZmZnd3d4iIiIiIiIiIiIiIiIiIiJmZmZmZmZmZmaqqqru7u93d3e7u7u7u7v///////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMy7u7vMzMy7u7u7u7u7u7u7u7uqqqqqqqqqqqqqqqqZmZmZmZmZmZmqqqqqqqq7u7u7u7u7u7uqqqqqqqqqqqqqqqq7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7vMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7uqqqq7u7u7u7u7u7vMzMzMzMzMzMzMzMzd3d3d3d3MzMzMzMzMzMzMzMzMzMy7u7vMzMy7u7u7u7u7u7uqqqqqqqqqqqp3d3dmZmZmZmZVVVVVVVVVVVVERERVVVVERERERERVVVV3d3dmZmZmZmZ3d3d3d3eIiIiIiIiIiIiZmZmIiIiZmZmZmZmIiIiIiIiIiIiIiIiIiIiIiIiZmZmZmZmZmZmZmZmZmZmIiIiZmZmIiIiIiIh3d3dmZmZmZmZVVVVVVVVERERERERERERERERERERERERERERERERERERVVVVVVVVERERERERVVVVmZmZ3d3d3d3eIiIiZmZmIiIiIiIiIiIiIiIiZmZmIiIiIiIh3d3dmZmZEREREREQzMzNERERERERVVVVmZmZmZmZVVVVVVVV3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIh3d3d3d3dmZmZmZmZmZmZERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZERERERERERERERERERERVVVVVVVVVVVVEREREREQzMzNERERERERERERmZmZ3d3eIiIiqqqrMzMzu7u7u7u7u7u7u7u7u7u7u7u7////u7u7u7u7u7u7////u7u7////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3MzMzMzMy7u7vMzMy7u7u7u7u7u7vMzMy7u7vMzMy7u7vMzMy7u7uqqqqIiIh3d3eIiIh3d3eIiIiZmZmIiIiZmZmIiIh3d3d3d3d3d3d3d3eIiIiIiIiZmZmqqqq7u7u7u7vd3d3d3d3u7u7d3d3d3d3d3d3d3d3u7u7d3d3d3d3MzMyqqqqIiIhmZmZmZmZEREREREQzMzMzMzMzMzNEREQzMzMzMzMzMzNEREQzMzNEREQzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzNEREQzMzNEREREREREREQzMzMiIiIzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzNERERmZmZmZmZVVVVVVVVmZmZmZmZmZmZ3d3dmZmZVVVVVVVVERERVVVVEREQzMzNERERERERVVVVVVVVVVVVmZmZ3d3dmZmZERERVVVVVVVVERERERERERERERERERERERERVVVVmZmZVVVVVVVVVVVVERERERERmZmZ3d3dmZmZVVVVVVVVVVVVVVVVEREREREQzMzNERERERERERERERERERERERERERERERERERERERERVVVV3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVUzMzNERERERERVVVVmZmZmZmZVVVVERERERERVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVmZmZmZmZmZmZVVVVERERERERERERVVVVVVVVVVVVVVVVEREREREQzMzNERERERERERERERERVVVVVVVVmZmZVVVVmZmZmZmaIiIiIiIhmZmZ3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZmIiIiIiIiIiIiIiIh3d3dmZmZVVVVVVVVERERERERmZmZ3d3eZmZmIiIiIiIh3d3eIiIh3d3d3d3d3d3dVVVVVVVVVVVVERERERERVVVVVVVVEREREREQzMzNEREQzMzMzMzNVVVV3d3dmZmZmZmZmZmZmZmZVVVVEREREREQzMzMzMzNERERERERERERERERERERERERERERERERERERVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3dmZmZmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVERERERERERERERERERERERERVVVVEREREREQzMzMzMzNEREQzMzMzMzMzMzNEREQzMzMzMzMzMzNERERVVVVVVVVVVVVERERERERERERERERVVVVVVVVEREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzNERERVVVVERERERERERERERERERERERERERERVVVVEREREREQzMzNEREQzMzNEREQzMzNERERERERERERERERERERERERVVVVVVVVVVVVVVVVERERVVVVERERERERERERVVVVVVVVERERVVVVEREQzMzMzMzMzMzNEREREREREREREREREREREREREREREREREREREREREREQzMzNEREQzMzNEREREREREREREREREREQzMzMzMzMiIiIiIiIzMzMzMzMzMzMiIiIzMzMiIiIzMzMiIiIzMzMzMzMzMzNERERERERVVVVVVVVVVVVERERERERVVVVVVVVVVVVERERERERERERERERERERERERERERERERERERERERERERERERERERVVVVVVVVEREQzMzNERERERERVVVVVVVVVVVVEREREREREREQzMzNEREQzMzNERERERERVVVVERERVVVVEREREREREREREREQzMzNERERVVVVmZmZVVVVmZmZmZmZVVVVERERVVVVmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVEREREREREREREREREREREREQzMzNVVVV3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVERERmZmZmZmZVVVVEREREREREREREREQzMzMiIiIzMzNEREREREQzMzMzMzMzMzMzMzMzMzNERERVVVVEREQzMzMzMzMzMzMzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzNEREREREQzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzNERERVVVVVVVVVVVUzMzNEREQzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREREREREREREREREREREREREREREREREREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzNERERmZmZVVVUzMzNEREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMiIiIiIiIREREzMzMzMzMiIiIzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzNERERVVVVVVVVmZmZ3d3dmZmZVVVV3d3d3d3d3d3eIiIh3d3eIiIiZmZmZmZmZmZmZmZmqqqrMzMzu7u7u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////7u7u7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzMzMzMzMzMu7u7u7u7u7u7zMzMzMzMzMzMzMzMu7u7qqqqu7u7u7u7qqqqu7u7u7u7u7u7qqqqqqqqqqqqqqqqu7u7u7u7qqqqu7u7qqqqmZmZqqqqqqqqu7u7u7u7u7u7u7u7zMzMzMzMu7u7zMzMzMzMzMzMzMzMzMzM3d3dzMzMzMzMzMzMzMzMzMzM3d3dzMzM3d3d3d3d3d3d3d3dzMzM3d3d3d3dzMzMzMzMzMzMu7u7u7u7qqqqu7u7qqqqu7u7u7u7u7u7u7u7u7u7zMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7qqqqmZmZiIiId3d3ZmZmZmZmZmZmVVVVVVVVREREVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmd3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiImZmZmZmZmZmZiIiIiIiImZmZiIiImZmZiIiIiIiIiIiId3d3d3d3d3d3ZmZmVVVVREREREREREREREREREREMzMzREREREREVVVVREREREREVVVVVVVVVVVVZmZmZmZmd3d3d3d3d3d3ZmZmd3d3iIiIiIiIiIiIiIiId3d3ZmZmREREREREREREZmZmVVVVZmZmVVVVREREREREd3d3d3d3d3d3ZmZmd3d3d3d3iIiId3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREREREVVVVZmZmZmZmZmZmVVVVVVVVREREREREMzMzVVVVVVVVVVVVVVVVVVVVREREREREREREMzMzMzMzREREVVVVd3d3mZmZu7u73d3d7u7u7u7u////7u7u////////7u7u////7u7u7u7u////7u7u7u7u////7u7u////////7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMu7u7zMzMu7u7qqqqmZmZqqqqmZmZmZmZiIiIiIiIiIiIiIiImZmZqqqqqqqqu7u7zMzMzMzMzMzM3d3dzMzMzMzMu7u7qqqqmZmZiIiImZmZmZmZqqqqiIiId3d3ZmZmVVVVREREMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREVVVVREREREREMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzREREREREREREIiIiMzMzMzMzREREVVVVZmZmZmZmVVVVZmZmVVVVVVVVZmZmZmZmREREVVVVVVVVVVVVREREREREREREREREREREREREVVVVVVVVd3d3ZmZmd3d3VVVVREREREREREREREREREREVVVVREREVVVVVVVVREREVVVVVVVVZmZmZmZmVVVVZmZmd3d3d3d3ZmZmVVVVVVVVREREREREVVVVVVVVVVVVVVVVREREVVVVREREREREREREREREREREVVVVVVVVZmZmZmZmZmZmVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmREREREREREREVVVVVVVVVVVVVVVVREREREREVVVVVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVREREVVVVZmZmZmZmVVVVVVVVVVVVREREVVVVREREREREREREVVVVVVVVVVVVZmZmVVVVZmZmZmZmd3d3d3d3VVVVd3d3d3d3iIiIiIiIiIiImZmZiIiIiIiIiIiImZmZmZmZmZmZiIiIiIiIiIiId3d3ZmZmVVVVVVVVMzMzMzMzZmZmd3d3mZmZiIiIiIiId3d3d3d3d3d3ZmZmZmZmZmZmVVVVVVVVVVVVREREREREREREREREMzMzREREREREREREREREREREd3d3d3d3d3d3ZmZmZmZmVVVVREREREREREREREREMzMzREREREREREREVVVVREREREREREREREREREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVREREVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREVVVVREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREVVVVZmZmREREREREMzMzREREVVVVREREVVVVREREREREVVVVMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzREREREREREREMzMzMzMzVVVVVVVVVVVVREREREREMzMzMzMzMzMzREREMzMzREREMzMzREREMzMzREREREREVVVVREREREREREREREREREREREREREREREREVVVVREREVVVVREREREREREREMzMzMzMzMzMzREREREREREREREREVVVVVVVVREREREREREREMzMzREREREREREREREREREREVVVVREREREREMzMzIiIiIiIiIiIiMzMzMzMzIiIiMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVREREVVVVZmZmVVVVZmZmVVVVVVVVREREREREREREREREREREREREREREMzMzREREREREMzMzREREVVVVVVVVREREMzMzMzMzVVVVVVVVVVVVZmZmVVVVREREREREREREMzMzREREREREREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVZmZmVVVVVVVVREREVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVREREREREMzMzMzMzREREZmZmd3d3ZmZmZmZmZmZmZmZmREREREREREREVVVVZmZmVVVVZmZmd3d3ZmZmVVVVd3d3d3d3REREMzMzREREMzMzIiIiMzMzMzMzMzMzMzMzREREMzMzMzMzREREREREREREREREREREMzMzMzMzIiIiIiIiMzMzIiIiREREVVVVMzMzMzMzMzMzMzMzMzMzREREREREMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVVVVVREREVVVVMzMzMzMzMzMzREREREREMzMzREREMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREREREMzMzREREMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREMzMzREREREREMzMzMzMzIiIiMzMzMzMzREREREREMzMzMzMzREREMzMzREREREREREREREREREREREREREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzREREREREZmZmVVVVREREREREVVVVREREREREMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzMzMzMzMzMzMzIiIiIiIiMzMzMzMzMzMzIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiERERIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREVVVVVVVVd3d3ZmZmZmZmZmZmd3d3ZmZmd3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiImZmZu7u73d3d7u7u7u7u7u7u////////////////7u7u////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////+7u7v///+7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3e7u7u7u7t3d3czMzN3d3czMzMzMzN3d3czMzMzMzMzMzLu7u8zMzLu7u7u7u7u7u6qqqru7u7u7u6qqqqqqqpmZmZmZmZmZmaqqqqqqqqqqqqqqqqqqqqqqqru7u7u7u7u7u8zMzMzMzMzMzMzMzN3d3d3d3czMzN3d3czMzMzMzN3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqru7u7u7u7u7u7u7u8zMzMzMzMzMzLu7u8zMzLu7u7u7u7u7u7u7u7u7u6qqqpmZmYiIiHd3d2ZmZmZmZlVVVVVVVVVVVVVVVWZmZlVVVVVVVWZmZlVVVVVVVWZmZnd3d2ZmZmZmZmZmZnd3d3d3d3d3d4iIiIiIiIiIiJmZmZmZmZmZmZmZmYiIiIiIiIiIiJmZmYiIiIiIiIiIiIiIiHd3d3d3d2ZmZmZmZlVVVVVVVURERERERERERDMzM0RERERERERERERERFVVVVVVVURERFVVVWZmZmZmZlVVVVVVVURERGZmZmZmZmZmZnd3d4iIiHd3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVURERERERHd3d3d3d1VVVWZmZmZmZnd3d3d3d3d3d3d3d2ZmZnd3d2ZmZnd3d4iIiHd3d3d3d2ZmZkRERERERERERFVVVVVVVWZmZlVVVWZmZmZmZmZmZlVVVURERERERFVVVVVVVWZmZlVVVVVVVURERFVVVURERERERDMzMzMzM0RERFVVVXd3d4iIiLu7u93d3e7u7v///////////////+7u7u7u7u7u7u7u7u7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u6qqqqqqqru7u7u7u8zMzMzMzN3d3czMzN3d3czMzMzMzLu7u6qqqpmZmXd3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVURERDMzMzMzMyIiIjMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIjMzMyIiIiIiIiIiIhERESIiIiIiIjMzMyIiIiIiIiIiIjMzMzMzM1VVVURERDMzMzMzM0RERERERDMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzM0RERERERDMzM0RERDMzMyIiIkRERERERERERDMzM0RERDMzMyIiIkRERDMzMzMzMzMzM0RERFVVVVVVVWZmZnd3d3d3d2ZmZmZmZlVVVWZmZkRERERERFVVVURERERERERERERERERERERERERERFVVVVVVVURERERERERERGZmZnd3d1VVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVWZmZlVVVURERGZmZoiIiGZmZlVVVVVVVVVVVURERFVVVVVVVWZmZlVVVURERFVVVURERFVVVURERERERERERERERERERFVVVWZmZlVVVVVVVVVVVVVVVWZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVURERERERFVVVWZmZlVVVURERERERERERERERERERERERERERFVVVURERFVVVURERFVVVWZmZlVVVVVVVVVVVURERFVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVURERFVVVWZmZmZmZnd3d1VVVVVVVWZmZlVVVVVVVWZmZmZmZnd3d4iIiIiIiIiIiJmZmZmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiIiIiHd3d2ZmZkRERERERDMzM0RERFVVVXd3d5mZmYiIiHd3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVURERFVVVVVVVTMzMzMzM0RERERERFVVVURERDMzM0RERGZmZnd3d3d3d3d3d1VVVVVVVVVVVURERERERERERERERERERFVVVVVVVURERERERFVVVURERERERERERFVVVVVVVVVVVWZmZmZmZnd3d2ZmZmZmZnd3d3d3d2ZmZmZmZlVVVVVVVVVVVWZmZlVVVVVVVWZmZlVVVVVVVURERFVVVVVVVWZmZlVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVURERDMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERDMzM1VVVVVVVVVVVURERERERERERERERFVVVURERERERERERERERDMzM0RERERERERERDMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVURERERERERERDMzMzMzMzMzM0RERDMzM0RERERERERERERERERERERERERERERERFVVVURERERERERERERERERERERERERERERERERERFVVVURERERERDMzMyIiIiIiIjMzM0RERERERERERERERERERERERERERERERDMzM0RERERERERERERERFVVVURERFVVVVVVVTMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzM0RERERERERERERERDMzM2ZmZnd3d3d3d2ZmZmZmZlVVVURERERERERERERERERERERERERERERERERERERERERERERERERERFVVVURERDMzM0RERERERFVVVWZmZmZmZlVVVVVVVURERERERERERDMzM0RERERERFVVVURERDMzM0RERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVURERERERERERDMzM0RERERERGZmZmZmZmZmZlVVVWZmZkRERERERERERERERFVVVWZmZlVVVXd3d3d3d4iIiGZmZmZmZmZmZjMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERERERDMzMyIiIjMzMyIiIhERESIiIiIiIiIiIiIiIkRERFVVVURERCIiIjMzMzMzMzMzM1VVVVVVVTMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzM0RERDMzM0RERERERERERERERDMzM0RERDMzM0RERDMzM0RERDMzMzMzMzMzM0RERDMzM0RERDMzM0RERERERDMzMzMzMyIiIjMzM0RERDMzM0RERERERERERDMzMzMzM0RERDMzMzMzM0RERERERDMzM0RERFVVVURERERERDMzMzMzM0RERDMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVVVVVURERERERERERERERDMzM0RERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERGZmZmZmZkRERERERFVVVURERDMzMzMzMzMzMzMzM0RERDMzM0RERDMzM0RERERERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIiIiIjMzMzMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERFVVVWZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d5mZmYiIiHd3d3d3d5mZmbu7u93d3f///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3u7u7d3d3d3d3d3d3MzMzd3d3MzMzd3d3d3d3d3d3d3d3u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3MzMzd3d3MzMzMzMzMzMzMzMzMzMzMzMzd3d3MzMzMzMzMzMy7u7u7u7uqqqqqqqqZmZmZmZmZmZmZmZmZmZmqqqqqqqqZmZmZmZmZmZmqqqqqqqqqqqqqqqqqqqqqqqqqqqq7u7vMzMy7u7vMzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3MzMzMzMzMzMzd3d3MzMy7u7vMzMzMzMzMzMy7u7u7u7vMzMy7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7uqqqq7u7u7u7uqqqqqqqq7u7uqqqqZmZmZmZmIiIiIiIhmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZ3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIh3d3eIiIh3d3d3d3d3d3dmZmZmZmZVVVVVVVVVVVVERERERERVVVVVVVVVVVVERERVVVVmZmZVVVVVVVVERERERERVVVVmZmZmZmZmZmZVVVVmZmZmZmZmZmZ3d3dmZmZ3d3d3d3dVVVVVVVUzMzNVVVV3d3dVVVUzMzNERER3d3dmZmZVVVVmZmZ3d3d3d3dmZmZ3d3d3d3d3d3dmZmZ3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVERERVVVUzMzNEREREREQiIiIzMzMzMzNERERERER3d3eZmZmqqqrd3d3u7u7u7u7////u7u7u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7d3d3d3d3MzMzMzMzMzMzMzMzMzMy7u7u7u7uqqqqZmZmZmZmqqqqqqqq7u7u7u7uqqqqZmZmIiIh3d3d3d3dmZmZmZmZVVVVERERERERVVVVEREREREREREQzMzMzMzMzMzMzMzMiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIiIiIzMzMzMzMiIiIiIiIiIiIzMzNEREQzMzMzMzMzMzNERERERERVVVVEREQzMzMzMzMiIiIzMzMiIiIzMzNERERERERERERVVVVEREREREREREQzMzNEREQzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzNERERERERERERVVVVVVVV3d3eIiIiIiIhmZmZ3d3dmZmZmZmZVVVVERERERERERERERERVVVVVVVVVVVVERERmZmZVVVVVVVVERERVVVV3d3d3d3d3d3dmZmZVVVVVVVVERERVVVVVVVVVVVVERERERERVVVVVVVVVVVVEREQzMzNERERVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZEREREREQzMzNVVVVmZmZVVVVVVVVmZmZVVVVmZmZ3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3dmZmZVVVVERERERERVVVVmZmZmZmZVVVVERERERERVVVVERERVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3dmZmZmZmZVVVVVVVVERERERERVVVVVVVV3d3eIiIiIiIiZmZmqqqqqqqqqqqqZmZmZmZmIiIiIiIiIiIiIiIiIiIh3d3dmZmZVVVVERERERERERERERERmZmaIiIiIiIh3d3eIiIh3d3d3d3d3d3dmZmZmZmZVVVVVVVVVVVVEREREREREREREREREREREREREREREREREREQzMzNERERVVVVmZmZmZmZmZmZVVVVERERERERVVVVERERERERVVVVVVVVVVVVERERERERERERERERERERERERERERERERVVVVVVVVmZmZmZmZ3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVERERERERERERVVVVVVVVmZmZVVVVmZmZVVVVVVVVVVVVEREREREQzMzNEREQzMzMzMzNERERERERVVVUzMzNEREQzMzMzMzMzMzNVVVVVVVVmZmZVVVVVVVVVVVVVVVVEREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVUzMzMzMzMzMzNERERERERVVVVVVVVEREREREREREREREQzMzNEREREREREREREREQzMzNERERERERERERERERERERERERERERERERERERVVVVERERERERERERERERVVVVVVVVVVVVEREREREREREQzMzMiIiIzMzMzMzMzMzMzMzNEREQzMzNEREQzMzNEREREREREREREREQzMzMzMzNERERERERERERVVVVVVVUzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzNEREREREQzMzMzMzNERERmZmZ3d3dmZmZVVVVVVVVVVVVVVVVERERERERERERERERERERERERERERERERERERERERVVVVVVVVEREQzMzNERERVVVVERERERERVVVVVVVVEREREREREREQzMzNEREREREREREREREREREREREREREREREREREREREREREQzMzNVVVVVVVVmZmZmZmZVVVVVVVVERERERERVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVVERERVVVVERERVVVVmZmZmZmZVVVVERERERERERERERERVVVVVVVVVVVVmZmZmZmZVVVVERERVVVVVVVVmZmZVVVVVVVVmZmZ3d3dmZmZVVVVVVVUzMzMzMzMzMzMzMzMzMzNERERVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIREREREREiIiIiIiIREREiIiIiIiIiIiJERERVVVUzMzMzMzMiIiIzMzMzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzNEREREREQzMzMzMzMiIiIzMzMzMzMzMzNERERVVVVVVVUzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzNEREQzMzNEREQzMzMzMzMzMzNERERERERERERERERVVVVVVVVEREREREREREQzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNVVVVmZmZVVVVEREREREREREQzMzNERERERERERERVVVVEREREREREREQzMzMzMzMzMzMzMzNERERERERmZmZVVVVVVVVERERERERERERERERERERVVVVVVVVERERERERERERERERVVVVERERERERERERERERVVVVEREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIzMzNEREQzMzNEREREREREREREREREREQzMzNERERVVVVmZmZmZmZVVVVERERVVVVVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIjMzMzu7u7////u7u7////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////7u7u3d3d3d3d3d3d3d3d3d3d7u7u3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzM3d3d3d3d3d3dzMzM3d3d3d3dzMzMzMzMzMzMzMzMu7u7u7u7qqqqqqqqqqqqqqqqmZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZmZmZmZmZmZmZmZmZu7u7qqqqu7u7u7u7u7u7u7u7zMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7zMzMzMzMzMzMu7u7zMzMu7u7u7u7u7u7qqqqu7u7qqqqqqqqqqqqqqqqqqqqqqqqqqqqu7u7qqqqqqqqqqqqqqqqqqqqqqqqiIiIiIiId3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVd3d3iIiIZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVd3d3d3d3ZmZmZmZmVVVVVVVVZmZmREREMzMzVVVVZmZmVVVVMzMzREREZmZmd3d3VVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmVVVVZmZmVVVVREREVVVVVVVVZmZmZmZmd3d3ZmZmVVVVVVVVVVVVREREREREMzMzREREREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzREREVVVVd3d3mZmZqqqqzMzMzMzM3d3d3d3d3d3d7u7u7u7u7u7u3d3d7u7u3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMu7u7zMzMzMzMzMzMu7u7qqqqmZmZiIiIiIiIiIiId3d3d3d3d3d3ZmZmZmZmd3d3ZmZmZmZmZmZmVVVVVVVVREREREREMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiERERIiIiERERERERERERIiIiIiIiIiIiIiIiIiIiIiIiMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREVVVVVVVVREREREREMzMzMzMzMzMzREREREREREREVVVVVVVVVVVVVVVVVVVVREREVVVVMzMzMzMzMzMzREREREREMzMzREREMzMzREREMzMzMzMzREREREREMzMzVVVVd3d3d3d3d3d3d3d3VVVVVVVVVVVVREREREREMzMzREREVVVVVVVVVVVVZmZmVVVVVVVVVVVVREREVVVVd3d3d3d3d3d3ZmZmVVVVVVVVVVVVREREREREVVVVVVVVVVVVREREREREVVVVREREMzMzMzMzREREVVVVVVVVREREREREREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVd3d3VVVVREREREREVVVVZmZmVVVVZmZmZmZmZmZmZmZmd3d3ZmZmd3d3d3d3iIiIiIiIiIiIiIiIZmZmVVVVVVVVREREVVVVZmZmd3d3ZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmVVVVZmZmd3d3ZmZmVVVVVVVVVVVVZmZmZmZmd3d3ZmZmd3d3d3d3d3d3ZmZmd3d3VVVVVVVVMzMzMzMzREREVVVVd3d3iIiImZmZqqqqmZmZmZmZqqqqqqqqqqqqmZmZiIiIiIiIiIiId3d3ZmZmZmZmREREREREREREVVVVVVVVVVVVZmZmd3d3iIiId3d3iIiId3d3ZmZmZmZmVVVVZmZmREREREREMzMzREREVVVVVVVVREREREREMzMzMzMzREREMzMzMzMzREREVVVVZmZmZmZmVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmREREREREREREMzMzREREREREREREREREVVVVVVVVVVVVVVVVZmZmZmZmd3d3VVVVVVVVd3d3ZmZmZmZmVVVVZmZmVVVVREREVVVVVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVREREMzMzMzMzVVVVZmZmZmZmVVVVZmZmZmZmREREREREREREREREREREMzMzREREMzMzREREVVVVVVVVREREREREMzMzMzMzIiIiREREVVVVZmZmZmZmZmZmZmZmREREREREMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzREREMzMzMzMzREREVVVVVVVVVVVVVVVVVVVVREREREREMzMzREREREREREREREREMzMzREREREREREREREREREREREREREREREREZmZmVVVVREREREREREREVVVVVVVVREREVVVVVVVVMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzMzMzREREMzMzMzMzMzMzREREMzMzMzMzIiIiMzMzMzMzREREREREVVVVMzMzMzMzIiIiMzMzMzMzIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVREREVVVVREREREREREREVVVVREREVVVVREREVVVVREREREREMzMzREREMzMzREREVVVVVVVVREREREREREREREREMzMzREREREREREREREREREREREREREREREREREREREREMzMzMzMzREREVVVVZmZmVVVVVVVVVVVVREREVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVREREREREVVVVVVVVZmZmVVVVREREREREREREREREVVVVVVVVVVVVd3d3ZmZmVVVVVVVVZmZmZmZmVVVVVVVVVVVVZmZmd3d3VVVVMzMzMzMzIiIiMzMzMzMzREREREREREREREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiERERIiIiERERERERIiIiERERIiIiIiIiERERREREVVVVMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzVVVVVVVVVVVVMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREVVVVZmZmVVVVREREREREMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREZmZmd3d3VVVVREREVVVVVVVVREREREREREREREREREREREREMzMzMzMzREREMzMzMzMzMzMzVVVVVVVVVVVVREREREREREREREREMzMzREREVVVVREREREREREREREREVVVVREREVVVVREREVVVVREREREREREREREREREREREREREREREREREREREREREREREREREREMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzMzMzMzMzMzMzIiIiREREREREVVVVZmZmVVVVREREVVVVREREREREREREVVVVVVVVZmZmVVVVREREREREVVVVZmZmZmZmd3d3ZmZmVVVVZmZmd3d3d3d3d3d3ZmZmVVVViIiIu7u73d3d////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////+7u7t3d3czMzN3d3d3d3d3d3czMzLu7u7u7u8zMzMzMzN3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3czMzN3d3czMzMzMzN3d3czMzN3d3czMzN3d3d3d3czMzMzMzN3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzN3d3czMzN3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzLu7u7u7u6qqqqqqqqqqqqqqqpmZmZmZmYiIiIiIiIiIiJmZmYiIiIiIiIiIiIiIiIiIiJmZmaqqqpmZmaqqqqqqqqqqqqqqqru7u7u7u6qqqru7u7u7u7u7u7u7u6qqqru7u8zMzMzMzLu7u8zMzMzMzLu7u7u7u7u7u7u7u6qqqru7u6qqqru7u6qqqpmZmZmZmaqqqpmZmaqqqpmZmaqqqqqqqqqqqpmZmZmZmZmZmYiIiIiIiHd3d3d3d2ZmZlVVVVVVVVVVVURERFVVVVVVVWZmZmZmZmZmZmZmZmZmZnd3d3d3d1VVVWZmZlVVVWZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVXd3d5mZmXd3d2ZmZlVVVWZmZmZmZlVVVURERERERFVVVWZmZlVVVWZmZmZmZlVVVVVVVVVVVVVVVURERFVVVURERDMzM0RERFVVVVVVVURERFVVVVVVVVVVVVVVVWZmZmZmZlVVVWZmZmZmZmZmZnd3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d1VVVVVVVVVVVURERDMzM0RERERERERERERERDMzMyIiIjMzMzMzMzMzMzMzM0RERDMzMzMzM0RERGZmZmZmZnd3d3d3d4iIiJmZmZmZmaqqqqqqqqqqqqqqqqqqqpmZmYiIiIiIiIiIiIiIiHd3d4iIiHd3d4iIiIiIiIiIiHd3d2ZmZlVVVVVVVURERERERFVVVVVVVURERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIhERERERERERERERERERESIiIiIiIhERERERESIiIhERESIiIiIiIiIiIhERESIiIhERERERESIiIhERESIiIiIiIiIiIiIiIhERESIiIjMzM0RERERERDMzMzMzMyIiIiIiIjMzMzMzMzMzMzMzM0RERERERDMzM0RERERERERERDMzM0RERERERERERFVVVVVVVWZmZlVVVVVVVVVVVVVVVURERERERDMzMyIiIkRERERERDMzM0RERDMzM0RERERERERERFVVVVVVVURERERERFVVVWZmZnd3d3d3d2ZmZlVVVVVVVURERERERERERERERERERFVVVVVVVVVVVVVVVURERERERERERERERFVVVURERFVVVURERERERERERERERERERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERFVVVVVVVURERFVVVVVVVVVVVWZmZlVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVURERERERFVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d4iIiIiIiHd3d4iIiIiIiHd3d2ZmZlVVVURERFVVVVVVVXd3d2ZmZlVVVVVVVWZmZlVVVVVVVWZmZmZmZmZmZnd3d3d3d2ZmZnd3d3d3d2ZmZmZmZmZmZnd3d3d3d3d3d2ZmZlVVVVVVVWZmZmZmZmZmZmZmZnd3d3d3d3d3d2ZmZnd3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZoiIiKqqqqqqqpmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiIiIiGZmZmZmZlVVVURERFVVVURERFVVVURERFVVVXd3d3d3d2ZmZnd3d4iIiHd3d1VVVVVVVWZmZlVVVVVVVURERERERERERFVVVVVVVURERDMzM0RERERERDMzMzMzMzMzM0RERERERFVVVVVVVVVVVVVVVURERFVVVVVVVWZmZmZmZmZmZlVVVVVVVURERERERERERERERDMzM0RERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVURERERERDMzMzMzM0RERGZmZlVVVWZmZmZmZlVVVVVVVVVVVVVVVTMzM0RERDMzM0RERDMzM0RERERERERERERERFVVVURERDMzMzMzMzMzM0RERHd3d2ZmZnd3d2ZmZlVVVURERERERDMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVVVVVVVVVWZmZlVVVVVVVTMzM0RERERERERERERERERERERERERERERERERERERERERERFVVVURERFVVVWZmZlVVVTMzM0RERERERERERERERFVVVVVVVURERERERDMzM0RERERERERERDMzMzMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMyIiIjMzMyIiIkRERFVVVTMzMzMzMyIiIjMzMyIiIjMzMyIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIkRERGZmZmZmZlVVVVVVVURERFVVVVVVVURERERERERERFVVVURERFVVVURERERERERERFVVVURERERERERERERERDMzM0RERERERERERFVVVVVVVURERDMzMzMzM0RERERERFVVVURERERERERERERERERERERERDMzM0RERDMzM0RERFVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVWZmZlVVVVVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVURERERERERERFVVVVVVVWZmZlVVVVVVVURERFVVVVVVVVVVVURERGZmZnd3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZjMzMzMzMzMzM0RERDMzM0RERERERERERERERDMzMzMzMzMzMyIiIjMzMzMzMyIiIiIiIiIiIhERERERESIiIhERESIiIhERESIiIiIiIhERESIiIjMzM0RERDMzMyIiIjMzMyIiIjMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzM1VVVVVVVVVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM0RERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVVVVVTMzM0RERERERDMzMzMzMzMzM0RERERERDMzM0RERDMzM0RERERERGZmZnd3d2ZmZlVVVURERFVVVVVVVVVVVURERFVVVURERERERERERERERERERERERDMzM0RERERERFVVVWZmZkRERERERERERDMzM0RERFVVVURERFVVVURERERERERERERERFVVVURERERERERERFVVVURERERERERERERERERERERERERERERERERERERERFVVVURERFVVVURERERERDMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMzMzMyIiIhERESIiIjMzMzMzMzMzMyIiIkRERFVVVWZmZmZmZmZmZlVVVVVVVURERERERERERFVVVVVVVVVVVURERERERERERFVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d4iIiHd3d2ZmZlVVVXd3d7u7u93d3e7u7v///+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////u7u7////u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3MzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3d3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3MzMzd3d3MzMzd3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3MzMzd3d3MzMzMzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7uqqqqqqqqqqqqZmZmZmZmZmZmIiIiZmZmZmZmZmZmZmZmZmZmqqqqqqqqZmZmqqqqqqqq7u7uqqqqqqqqqqqqZmZmqqqq7u7uqqqq7u7u7u7u7u7u7u7u7u7u7u7uqqqq7u7uqqqq7u7u7u7uqqqqqqqqqqqqqqqqqqqqZmZmqqqqqqqqZmZmqqqqZmZmZmZmZmZmIiIiZmZmIiIiIiIiIiIh3d3d3d3dmZmZmZmZVVVVVVVVmZmZVVVVVVVVVVVVmZmZ3d3dmZmZmZmZ3d3dmZmZVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3d3d3d3d3eIiIh3d3d3d3d3d3dmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZ3d3d3d3d3d3d3d3d3d3dmZmZVVVVEREREREREREQzMzNERERVVVVmZmZmZmZVVVVmZmZmZmZmZmZVVVVVVVUzMzMzMzNEREREREQzMzNERERVVVVERERVVVVmZmZmZmZVVVVVVVVVVVV3d3d3d3d3d3dmZmZVVVVVVVVmZmZVVVVERERVVVVmZmZVVVVVVVVVVVVmZmZmZmZEREREREREREREREQzMzMzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNERERERERERERERERERERVVVVVVVVVVVVVVVVEREQzMzNERERERERERERVVVVERERERERERERERERVVVVEREREREQzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIREREREREiIiIiIiIREREREREiIiIREREiIiIiIiIREREREREREREREREiIiIREREREREiIiIREREiIiIREREiIiIREREREREREREREREiIiIREREiIiIiIiIiIiIiIiIREREREREiIiIREREREREiIiIiIiIREREiIiIiIiIiIiIiIiJEREREREREREQzMzMzMzNEREQzMzNERERERERVVVVEREREREREREQzMzNEREREREQzMzNEREREREREREQzMzMzMzNERERVVVVmZmZmZmZVVVVEREREREREREQzMzNEREQzMzMzMzMzMzMzMzNERERERERERERVVVVVVVVERERVVVVVVVVERERERERmZmaIiIh3d3dmZmZmZmZVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZERERVVVVEREQzMzMzMzNERERVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVERERERERERERERERVVVVVVVVERERVVVVVVVVVVVVmZmZVVVVVVVVmZmZ3d3dmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3eIiIiZmZmIiIiIiIiIiIiZmZlmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3dVVVVVVVVmZmZ3d3d3d3dmZmZmAP//AABmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZlVVVVVVVVVVVURERFVVVWZmZmZmZnd3d3d3d4iIiIiIiIiIiIiIiJmZmZmZmZmZmYiIiHd3d3d3d2ZmZmZmZmZmZlVVVURERFVVVVVVVURERERERFVVVWZmZoiIiIiIiHd3d3d3d4iIiGZmZlVVVVVVVVVVVURERFVVVVVVVVVVVWZmZlVVVURERERERERERDMzM0RERERERERERERERERERERERFVVVWZmZmZmZmZmZlVVVWZmZmZmZnd3d2ZmZlVVVURERERERDMzM0RERDMzM0RERERERERERFVVVVVVVVVVVVVVVVVVVURERFVVVWZmZnd3d2ZmZmZmZmZmZmZmZlVVVWZmZlVVVURERFVVVURERERERFVVVVVVVVVVVVVVVWZmZlVVVVVVVURERDMzM0RERERERFVVVVVVVXd3d2ZmZlVVVVVVVWZmZkRERERERERERERERDMzM0RERDMzMzMzM0RERFVVVVVVVWZmZkRERDMzMzMzM0RERFVVVXd3d3d3d2ZmZkRERDMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzM1VVVVVVVURERFVVVWZmZlVVVVVVVURERERERDMzM0RERDMzM0RERERERERERDMzM0RERERERFVVVURERFVVVURERFVVVVVVVTMzM0RERERERFVVVVVVVVVVVURERERERERERERERERERDMzMzMzM0RERDMzMyIiIjMzMyIiIjMzMzMzMyIiIjMzMzMzM1VVVURERDMzMyIiIiIiIjMzMzMzM1VVVTMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzM0RERDMzM0RERGZmZlVVVVVVVURERFVVVVVVVURERERERFVVVURERFVVVVVVVVVVVVVVVURERFVVVURERFVVVURERERERERERDMzM0RERFVVVVVVVVVVVURERFVVVURERERERERERFVVVVVVVVVVVURERERERERERERERDMzM0RERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVWZmZlVVVVVVVWZmZmZmZlVVVVVVVWZmZlVVVVVVVURERERERFVVVURERFVVVVVVVURERERERERERERERFVVVWZmZnd3d2ZmZnd3d2ZmZlVVVURERFVVVVVVVVVVVWZmZmZmZkRERDMzM0RERERERDMzM0RERERERERERDMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIhERERERERERESIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzM0RERERERDMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzM0RERGZmZlVVVTMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERERERDMzMyIiIjMzMzMzM0RERDMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzM0RERERERERERFVVVVVVVURERERERDMzM0RERERERDMzMzMzM0RERDMzM0RERDMzM0RERERERFVVVXd3d3d3d2ZmZlVVVURERFVVVURERFVVVVVVVURERFVVVVVVVURERERERERERDMzM0RERERERFVVVWZmZlVVVURERERERERERERERFVVVURERFVVVURERERERERERERERERERERERFVVVURERFVVVURERERERFVVVURERERERERERERERERERERERERERERERERERERERFVVVURERFVVVVVVVURERDMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIkRERGZmZmZmZmZmZmZmZlVVVURERFVVVURERFVVVVVVVVVVVURERERERERERERERFVVVWZmZlVVVWZmZmZmZmZmZmZmZnd3d3d3d3d3d2ZmZmZmZoiIiKqqqt3d3e7u7v///+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////u7u7u7u7d3d3u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3u7u7d3d3u7u7d3d3u7u7d3d3d3d3d3d3MzMzMzMzd3d3d3d3d3d3d3d3MzMzMzMzd3d3MzMzd3d3d3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMy7u7vMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3MzMzd3d3MzMzd3d3MzMzMzMzd3d3MzMzMzMy7u7uqqqqqqqqqqqqqqqqqqqqqqqqqqqqZmZmqqqqZmZmqqqqqqqqqqqqqqqqqqqqqqqqZmZmZmZmZmZmZmZmZmZmIiIiIiIiIiIiIiIiZmZmIiIiZmZmZmZmqqqqqqqqqqqqqqqq7u7u7u7uqqqq7u7uqqqq7u7uqqqqZmZmqqqqZmZmIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3eIiIiIiIh3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3eZmZmIiIh3d3dmZmZVVVVmZmZVVVVERERVVVVmZmZmZmZmZmZERERERERmZmZmZmZVVVVmZmZVVVVVVVUzMzMzMzMzMzMzMzMzMzMzMzNVVVWIiIh3d3dmZmZVVVVVVVVVVVVmZmZVVVVmZmZmZmZ3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVUzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIREREREREREREREREREREiIiIREREREREiIiIREREREREiIiIREREiIiIiIiIiIiIREREiIiIREREREREiIiIREREREREiIiIiIiIiIiIREREiIiIREREiIiIREREREREREREiIiIzMzMzMzMiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIzMzMiIiJEREREREQzMzNERERERERERERVVVVVVVVmZmZmZmZEREREREREREREREREREREREQzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzNVVVVmZmZmZmZmZmZVVVVVVVVERERVVVVEREQzMzNEREQzMzNERERERERERERVVVVERERERERERERVVVVVVVVERERERERVVVVVVVVmZmZmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dVVVVVVVVVVVVERERERERVVVVmZmZVVVVVVVVVVVVVVVVERERERERVVVVmZmZmZmZVVVVmZmZVVVVVVVUzMzNERERVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZ3d3d3d3dmZmZVVVVERERERERmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIiZmZmZmZmZmZmZmZmZmZmZmZmIiIiIiIhmZmZmZmZmZmZ3d3dmZmZmZmZVVVVmZmZmZmZ3d3d3d3d3d3dVVVVmZmZmZmZVVVVmZmZmZmZ3d3d3d3dmZmZVVVVVVVVmZmZ3d3eIiIiIiIh3d3d3d3d3d3d3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVERERERERmZmZmZmZmZmZmZmaIiIiIiIiIiIiIiIiZmZmZmZmIiIh3d3dVVVV3d3d3d3dmZmZmZmZVVVVmZmZVVVVVVVVERERVVVVVVVVVVVVmZmaIiIiIiIh3d3d3d3eIiIh3d3dmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVEREREREQzMzNEREQzMzNEREREREQzMzMzMzMzMzMzMzNmZmZmZmZ3d3dmZmZmZmZmZmZmZmZEREREREQzMzNEREQzMzNEREQzMzNERERERERERERVVVVVVVVVVVVVVVVVVVVERERERERVVVVmZmZ3d3d3d3dmZmZVVVVVVVVmZmZmZmZVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVmZmZVVVVVVVUzMzNERERVVVVERERVVVVmZmZVVVVVVVVmZmZVVVVVVVVEREREREREREQzMzNEREQzMzNERERERERVVVVVVVVmZmZVVVUzMzMzMzNERERmZmZ3d3dmZmZVVVVEREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERERERERERERERERERERERERERVVVVVVVVERERVVVVEREREREQzMzNERERVVVVERERVVVVEREQzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzNEREREREQzMzMzMzMzMzMiIiIiIiJEREREREQzMzMiIiIiIiIiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNVVVVVVVVVVVVVVVVERERERERVVVVERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVERERVVVVERERERERERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERERERERERERERVVVVERERERERERERERERVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZVVVVVVVVERERERERERERERERVVVVVVVVVVVVERERERERERERERERVVVV3d3eIiIiIiIhmZmZ3d3dmZmZmZmZVVVVVVVVVVVVEREREREREREREREREREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMiIiIREREREREREREREREiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIREREiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNVVVVVVVUzMzMzMzMzMzMzMzMiIiIzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERVVVVVVVVVVVVEREREREREREQzMzNEREREREREREREREREREREREREREQzMzNERER3d3d3d3d3d3d3d3dVVVVVVVVERERVVVVERERVVVVVVVVERERVVVVVVVVERERERERERERERERERERmZmZVVVVEREQzMzMzMzNERERVVVVVVVVEREREREQzMzNERERERERERERVVVVERERERERVVVVVVVVERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERVVVVVVVVEREREREQzMzMzMzMzMzMiIiIzMzMiIiIzMzNEREQiIiIREREiIiIiIiIiIiIzMzNERERmZmZ3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZmZmZVVVVVVVV3d3dmZmZERERVVVVmZmZ3d3d3d3d3d3dmZmZmZmZ3d3eIiIiqqqrMzMzu7u7u7u7////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMu7u7zMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7zMzMu7u7u7u7u7u7u7u7zMzMzMzMzMzMzMzMu7u7zMzMu7u7u7u7zMzMu7u7zMzMu7u7u7u7u7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqqqqqqqqqmZmZmZmZqqqqmZmZiIiIiIiId3d3ZmZmZmZmZmZmVVVVZmZmZmZmZmZmd3d3d3d3iIiIiIiImZmZmZmZmZmZqqqqqqqqqqqqqqqqqqqqqqqqqqqqmZmZiIiImZmZiIiIiIiIiIiId3d3iIiIiIiIiIiId3d3iIiId3d3iIiId3d3d3d3d3d3ZmZmZmZmZmZmVVVVREREVVVVREREVVVVVVVVREREVVVVZmZmVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmd3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3iIiIZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmVVVVREREREREVVVVREREVVVVVVVVVVVVREREVVVVREREREREREREMzMzMzMzVVVVd3d3d3d3d3d3VVVVREREREREVVVVVVVVVVVVZmZmZmZmd3d3VVVVVVVVVVVVZmZmREREREREREREREREREREREREVVVVZmZmZmZmMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiIiIiMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzMzMzMzMzIiIiIiIiERERIiIiERERERERIiIiERERIiIiERERIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiERERIiIiIiIiERERIiIiERERERERIiIiIiIiERERIiIiERERIiIiERERIiIiERERIiIiERERIiIiMzMzREREMzMzIiIiIiIiERERERERIiIiERERIiIiMzMzREREMzMzIiIiERERERERERERIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzREREVVVVVVVVZmZmZmZmiIiIZmZmREREVVVVVVVVREREMzMzMzMzMzMzREREREREMzMzMzMzMzMzREREMzMzREREREREZmZmd3d3d3d3d3d3VVVVVVVVREREMzMzMzMzMzMzMzMzREREVVVVVVVVVVVVREREREREVVVVVVVVVVVVREREVVVVZmZmZmZmZmZmVVVVVVVVZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVREREREREVVVVZmZmVVVVVVVVREREVVVVREREVVVVVVVVZmZmZmZmVVVVVVVVZmZmREREMzMzREREZmZmd3d3VVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmVVVVVVVVVVVVVVVVd3d3d3d3iIiIiIiIiIiId3d3d3d3iIiImZmZmZmZmZmZmZmZiIiIiIiIiIiId3d3d3d3ZmZmZmZmd3d3d3d3ZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmd3d3d3d3iIiIZmZmZmZmZmZmd3d3iIiIiIiId3d3d3d3d3d3d3d3ZmZmd3d3ZmZmZmZmZmZmd3d3ZmZmVVVVREREREREREREZmZmVVVVVVVVZmZmd3d3mZmZmZmZmZmZmZmZmZmZd3d3ZmZmZmZmZmZmd3d3ZmZmVVVVZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVViIiIiIiId3d3iIiId3d3ZmZmVVVVZmZmZmZmVVVVVVVVVVVVREREREREREREMzMzREREMzMzREREREREMzMzMzMzMzMzMzMzREREVVVViIiId3d3ZmZmd3d3ZmZmVVVVREREVVVVMzMzREREMzMzREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREd3d3d3d3d3d3ZmZmVVVVVVVVZmZmVVVVVVVVVVVVVVVVREREVVVVREREVVVVVVVVVVVVZmZmVVVVREREREREREREVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVREREREREREREREREREREMzMzMzMzREREREREVVVVVVVVVVVVVVVVMzMzREREZmZmZmZmZmZmVVVVVVVVREREREREREREREREREREMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREMzMzMzMzMzMzIiIiMzMzREREREREREREREREREREREREVVVVVVVVREREREREMzMzMzMzREREMzMzREREREREVVVVREREVVVVVVVVVVVVVVVVREREREREREREVVVVVVVVREREREREREREREREREREREREREREMzMzREREMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzREREMzMzIiIiMzMzIiIiMzMzMzMzVVVVMzMzIiIiIiIiERERERERIiIiERERIiIiERERIiIiIiIiMzMzIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzVVVVZmZmVVVVVVVVREREREREVVVVREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVREREREREMzMzREREREREREREREREVVVVVVVVVVVVVVVVREREREREREREVVVVVVVVZmZmZmZmVVVVVVVVVVVVREREVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVREREVVVVVVVVZmZmVVVVREREMzMzREREVVVVREREZmZmiIiImZmZVVVVZmZmiIiId3d3VVVVREREREREMzMzMzMzREREVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiERERIiIiERERERERIiIiERERERERIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzREREVVVVREREMzMzIiIiMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREMzMzREREMzMzMzMzREREREREREREVVVVVVVVREREVVVVREREREREMzMzREREMzMzREREREREREREREREREREREREVVVVd3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVVVVVVVVVREREMzMzMzMzREREVVVVVVVVVVVVREREREREREREREREREREREREREREREREREREREREREREVVVVREREREREREREREREREREREREREREREREREREREREREREREREVVVVREREREREREREREREREREREREREREMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzIiIiMzMzZmZmiIiId3d3d3d3VVVVZmZmVVVVVVVVd3d3iIiIiIiIZmZmd3d3d3d3ZmZmZmZmZmZmd3d3VVVVVVVVZmZmd3d3d3d3d3d3d3d3ZmZmd3d3iIiIiIiIqqqq3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////+7u7u7u7t3d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzN3d3czMzMzMzMzMzN3d3czMzMzMzMzMzMzMzMzMzLu7u8zMzMzMzMzMzN3d3d3d3czMzMzMzN3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u7u7u8zMzLu7u7u7u6qqqru7u6qqqru7u7u7u6qqqru7u6qqqqqqqqqqqqqqqru7u7u7u8zMzLu7u8zMzMzMzMzMzMzMzLu7u8zMzLu7u7u7u7u7u7u7u6qqqqqqqqqqqqqqqpmZmYiIiHd3d2ZmZlVVVVVVVVVVVURERERERERERFVVVVVVVVVVVVVVVWZmZmZmZnd3d3d3d3d3d3d3d4iIiIiIiIiIiJmZmZmZmZmZmZmZmZmZmYiIiIiIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiHd3d4iIiIiIiHd3d3d3d3d3d2ZmZmZmZlVVVVVVVURERFVVVURERERERFVVVURERFVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZnd3d2ZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZnd3d2ZmZnd3d3d3d4iIiIiIiHd3d3d3d2ZmZnd3d3d3d2ZmZlVVVWZmZkRERFVVVVVVVURERERERFVVVVVVVURERERERERERFVVVVVVVURERDMzM0RERFVVVXd3d2ZmZkRERDMzM0RERERERERERFVVVVVVVWZmZlVVVVVVVVVVVWZmZlVVVVVVVTMzM0RERERERERERERERFVVVVVVVVVVVURERERERERERERERCIiIjMzMzMzMzMzMyIiIiIiIjMzMzMzMyIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIhERESIiIhERERERESIiIhERESIiIhERERERERERERERESIiIiIiIhERESIiIhERERERESIiIhERESIiIiIiIhERESIiIhERERERESIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIhERERERERERESIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIhERESIiIhERESIiIiIiIjMzMzMzMzMzMyIiIhERESIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMyIiIjMzM0RERFVVVVVVVVVVVWZmZnd3d3d3d2ZmZlVVVVVVVVVVVTMzMzMzMzMzMzMzM0RERERERDMzMzMzMzMzM0RERDMzM0RERFVVVVVVVVVVVXd3d3d3d2ZmZkRERERERDMzMzMzMzMzMyIiIkRERFVVVVVVVVVVVURERERERFVVVURERERERERERFVVVVVVVWZmZmZmZlVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVVVVVURERERERFVVVWZmZlVVVVVVVURERFVVVVVVVWZmZnd3d3d3d2ZmZmZmZmZmZmZmZkRERERERERERGZmZnd3d2ZmZlVVVVVVVVVVVWZmZnd3d3d3d2ZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d4iIiIiIiIiIiHd3d3d3d4iIiIiIiJmZmZmZmZmZmYiIiIiIiIiIiIiIiHd3d2ZmZmZmZnd3d3d3d4iIiHd3d3d3d3d3d3d3d2ZmZoiIiHd3d3d3d3d3d2ZmZmZmZnd3d3d3d2ZmZmZmZmZmZlVVVWZmZoiIiIiIiHd3d3d3d4iIiHd3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVURERFVVVURERFVVVVVVVVVVVWZmZoiIiJmZmYiIiJmZmYiIiHd3d2ZmZmZmZmZmZnd3d2ZmZmZmZlVVVVVVVURERFVVVVVVVVVVVWZmZmZmZlVVVVVVVWZmZnd3d4iIiIiIiIiIiGZmZmZmZnd3d2ZmZkRERERERERERERERDMzM1VVVURERERERERERERERERERERERERERERERDMzMzMzM0RERHd3d3d3d3d3d2ZmZmZmZkRERFVVVVVVVURERERERERERERERERERERERERERERERFVVVVVVVVVVVVVVVURERDMzM1VVVWZmZnd3d2ZmZmZmZlVVVWZmZmZmZlVVVWZmZmZmZmZmZlVVVURERFVVVVVVVWZmZmZmZlVVVVVVVURERERERERERFVVVWZmZlVVVWZmZlVVVVVVVVVVVURERERERERERERERERERDMzMzMzMzMzMzMzM1VVVURERERERERERGZmZkRERERERHd3d2ZmZmZmZlVVVVVVVVVVVURERERERERERERERERERERERDMzM0RERDMzMzMzM0RERDMzM0RERDMzMyIiIjMzMzMzMzMzM0RERERERFVVVURERERERERERERERFVVVURERERERDMzM0RERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVURERERERERERFVVVURERFVVVURERERERDMzM0RERERERDMzMzMzMzMzM0RERERERDMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMyIiIjMzMyIiIjMzM0RERDMzMyIiIiIiIiIiIhERERERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzM0RERGZmZlVVVVVVVURERFVVVVVVVURERERERFVVVURERERERERERFVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVURERFVVVURERERERERERERERERERERERERERERERERERFVVVVVVVVVVVURERFVVVTMzM0RERERERGZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVURERFVVVVVVVURERERERERERERERERERERERFVVVWZmZlVVVTMzMzMzM0RERFVVVURERERERIiIiIiIiGZmZlVVVWZmZmZmZnd3d1VVVURERCIiIkRERFVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIhERESIiIhERERERESIiIhERESIiIhERERERESIiIiIiIjMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzM0RERERERERERDMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERERERERERDMzMzMzMyIiIjMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzM0RERERERERERERERFVVVURERFVVVURERDMzM0RERDMzM0RERERERERERERERERERERERGZmZnd3d2ZmZnd3d2ZmZmZmZlVVVWZmZlVVVURERFVVVWZmZlVVVWZmZlVVVVVVVVVVVURERERERFVVVWZmZlVVVTMzMzMzMzMzM1VVVWZmZlVVVURERERERERERDMzM0RERERERERERERERERERFVVVURERERERFVVVURERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERDMzMyIiIjMzMyIiIjMzMzMzMzMzMyIiIiIiIiIiIjMzMzMzM1VVVYiIiIiIiIiIiGZmZmZmZlVVVXd3d5mZmaqqqqqqqpmZmYiIiHd3d1VVVWZmZmZmZmZmZmZmZlVVVWZmZmZmZnd3d3d3d3d3d3d3d3d3d4iIiJmZmYiIiKqqqszMzN3d3e7u7v///////////////+7u7v///////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////u7u7////////////////////u7u7u7u7d3d3u7u7d3d3u7u7d3d3u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzd3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMy7u7uqqqq7u7u7u7u7u7u7u7vMzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7vMzMy7u7u7u7u7u7vMzMy7u7u7u7u7u7u7u7u7u7u7u7vMzMzMzMy7u7vMzMy7u7u7u7uqqqq7u7uqqqqqqqqqqqqZmZmqqqqqqqqqqqqqqqq7u7uqqqq7u7u7u7u7u7vMzMzMzMy7u7vMzMzMzMy7u7u7u7vMzMy7u7uqqqqqqqqZmZmIiIiIiIh3d3dmZmZVVVVVVVVERERERERERERERERERERERERERERERERVVVVERERVVVVVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3eIiIiIiIh3d3eIiIiIiIiIiIiIiIiIiIiZmZmIiIiIiIiIiIiIiIh3d3eIiIiIiIiIiIiIiIiIiIh3d3d3d3dmZmZmZmZmZmZVVVVVVVVVVVVVVVVERERERERERERVVVVVVVVmZmZVVVVVVVVmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3dmZmZmZmZmZmZ3d3d3d3dmZmZmZmZmZmZmZmZ3d3eIiIiIiIh3d3eIiIiZmZmIiIhmZmZ3d3eIiIiIiIhmZmZEREREREREREQzMzMzMzNERERVVVVEREQzMzNERERERERERERERERERERVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzNERERVVVVVVVVERERERERVVVVVVVVERERVVVVERERVVVVVVVVEREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIREREREREiIiIREREiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIREREiIiIREREREREiIiIREREiIiIiIiIREREiIiIiIiIzMzMzMzMiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIREREREREiIiIREREiIiIzMzNVVVVVVVUzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNERERVVVVVVVVVVVVVVVV3d3eIiIiIiIhmZmZERERVVVVmZmZVVVVEREREREQzMzMzMzNERERERERERERERERERERERERERERVVVVVVVVEREQzMzNVVVVEREREREREREREREQzMzMzMzNERERERERERERERERERERERERVVVVEREREREREREQzMzNERERERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZ3d3dmZmZmZmZmZmZmZmZVVVVERERERERVVVVVVVVmZmZVVVVVVVVmZmZVVVVVVVV3d3d3d3dmZmZ3d3d3d3d3d3d3d3dVVVVERERVVVV3d3eIiIh3d3dmZmZmZmZ3d3d3d3d3d3eIiIh3d3d3d3dmZmZmZmZVVVVmZmZVVVVmZmZ3d3d3d3eIiIiIiIiIiIiZmZmIiIiIiIiIiIiZmZmZmZmqqqqZmZmIiIiZmZmIiIiIiIh3d3dmZmZmZmZ3d3eIiIiZmZmIiIiZmZmIiIh3d3eIiIiIiIiIiIh3d3d3d3dmZmZmZmZmZmZmZmZVVVVVVVVERERVVVVERERmZmaIiIiIiIiIiIh3d3d3d3d3d3d3d3eIiIiIiIhmZmZ3d3d3d3d3d3dVVVVVVVVVVVVVVVVERERERERVVVVVVVVVVVVmZmaIiIiIiIiIiIiIiIiZmZl3d3d3d3dmZmZ3d3dmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVmZmaIiIh3d3d3d3dmZmZ3d3dmZmZVVVUzMzMzMzNERERERERERERERERERERERERERERVVVVEREQzMzNERERERERERERERERmZmaIiIh3d3dmZmZERERVVVVERERVVVVVVVVVVVVVVVVERERERERERERERERERERmZmZVVVVVVVVVVVVEREQzMzNVVVWIiIh3d3d3d3dmZmZVVVVmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVERERERERERERERERVVVVEREQzMzMzMzNEREQzMzMzMzNERERERERERERERERERERVVVVERERVVVVmZmZVVVVmZmZVVVVEREREREREREREREQzMzNEREREREREREREREREREREREREREQzMzMzMzMzMzMzMzNEREQzMzNERERERERERERVVVVEREREREQzMzNERERVVVVERERERERERERERERERERERERERERERERmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVEREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzNVVVVmZmZVVVVVVVVVVVVVVVVmZmZVVVVERERERERERERERERVVVVERERmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERmZmZVVVVVVVVERERVVVVERERERERERERERERERERERERERERERERVVVVERERVVVVERERERERERERERERERERERERmZmZVVVVVVVVVVVVVVVVERERERERERERERERERERERERERERVVVVVVVVERERERERERERERERERERERERERERERERVVVVERERERERERERVVVVEREQzMzNERERERERERERmZmZ3d3d3d3d3d3eIiIh3d3dmZmZEREQzMzNERERVVVVEREQzMzMzMzMzMzMzMzNERERVVVVEREQiIiIzMzNEREQzMzMiIiIREREiIiIREREiIiIREREREREREREiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMzMzNEREQzMzMzMzMzMzNVVVVEREQzMzMiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzNEREQzMzNEREREREREREQzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzNEREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzNERERmZmZVVVVEREREREREREREREREREQzMzNEREQzMzMzMzMzMzNERERVVVVERERmZmZ3d3dmZmZ3d3d3d3dVVVVVVVVVVVVVVVVERERmZmZmZmZ3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVmZmZEREQzMzNERERVVVVVVVVVVVVERERERERERERERERERERERERERERERERERERVVVVERERERERVVVVEREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREQzMzMzMzNEREREREQiIiIiIiIiIiIiIiIzMzMzMzNERERmZmaZmZmIiIiIiIhmZmZmZmZ3d3eZmZmqqqq7u7uZmZmZmZmIiIh3d3dVVVVVVVV3d3dmZmZVVVVmZmZmZmZmZmZmZmZ3d3eIiIh3d3d3d3d3d3eIiIiqqqqqqqqqqqq7u7vd3d3u7u7////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d3d3d7u7u3d3d7u7u7u7u7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqu7u7u7u7u7u7u7u7qqqqu7u7u7u7u7u7u7u7u7u7zMzMu7u7zMzMu7u7u7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqmZmZqqqqu7u7qqqqu7u7u7u7u7u7zMzMu7u7u7u7zMzMu7u7qqqqqqqqqqqqu7u7mZmZmZmZmZmZd3d3d3d3ZmZmZmZmVVVVVVVVVVVVREREREREREREREREREREREREREREREREREREREREVVVVREREVVVVVVVVZmZmZmZmVVVVZmZmd3d3ZmZmd3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZiIiImZmZiIiIiIiIiIiIiIiIiIiId3d3d3d3ZmZmZmZmZmZmZmZmVVVVVVVVREREVVVVREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3iIiIZmZmZmZmVVVVZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3iIiIiIiIiIiId3d3d3d3iIiImZmZd3d3VVVVVVVVVVVVMzMzMzMzZmZmZmZmREREMzMzREREREREMzMzREREREREREREMzMzREREREREMzMzMzMzIiIiMzMzREREREREMzMzMzMzREREREREREREREREVVVVVVVVVVVVREREREREVVVVVVVVREREREREREREREREREREMzMzMzMzIiIiMzMzREREREREIiIiMzMzREREREREMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzMzMzIiIiERERIiIiERERIiIiIiIiIiIiERERERERIiIiERERIiIiIiIiMzMzIiIiIiIiERERIiIiIiIiIiIiERERIiIiIiIiERERIiIiIiIiMzMzMzMzMzMzIiIiMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiERERERERIiIiERERERERERERMzMzVVVVZmZmVVVVREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVZmZmVVVVZmZmZmZmiIiIiIiIiIiIZmZmZmZmZmZmVVVVREREREREREREREREREREVVVVREREREREREREVVVVREREMzMzREREREREMzMzMzMzVVVVREREREREREREMzMzMzMzREREREREREREREREREREREREREREVVVVREREREREMzMzMzMzREREVVVVZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmREREVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmd3d3d3d3ZmZmZmZmZmZmVVVVVVVVd3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3iIiId3d3d3d3ZmZmZmZmZmZmZmZmVVVVREREd3d3mZmZiIiImZmZmZmZiIiIiIiIiIiImZmZmZmZqqqqqqqqmZmZmZmZmZmZiIiIiIiId3d3ZmZmVVVVd3d3iIiImZmZiIiIiIiIiIiIiIiId3d3d3d3d3d3iIiIiIiId3d3VVVVVVVVZmZmVVVVREREREREREREVVVVVVVVZmZmmZmZiIiId3d3d3d3iIiIiIiIiIiId3d3d3d3d3d3iIiIZmZmZmZmVVVVZmZmREREVVVVREREREREVVVVZmZmVVVVd3d3ZmZmd3d3iIiIiIiIiIiIZmZmZmZmd3d3ZmZmZmZmZmZmVVVVREREVVVVVVVVZmZmZmZmd3d3d3d3d3d3ZmZmREREREREVVVVd3d3d3d3iIiIiIiId3d3ZmZmVVVVREREREREMzMzREREREREREREMzMzREREREREREREVVVVREREREREMzMzMzMzVVVVZmZmd3d3d3d3VVVVVVVVREREVVVVREREVVVVVVVVREREREREREREREREREREVVVVVVVVVVVVVVVVREREREREREREVVVVd3d3d3d3d3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVZmZmVVVVZmZmZmZmZmZmREREMzMzVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREVVVVREREREREREREREREREREMzMzREREREREMzMzVVVVVVVVVVVVVVVVVVVVVVVVZmZmREREREREREREREREMzMzREREVVVVREREREREREREMzMzREREMzMzREREMzMzMzMzMzMzMzMzMzMzREREVVVVREREVVVVVVVVREREREREVVVVREREREREREREMzMzREREVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmREREREREREREMzMzREREREREMzMzMzMzMzMzMzMzREREREREREREREREMzMzMzMzMzMzREREMzMzMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiERERERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzVVVVZmZmZmZmVVVVVVVVVVVVREREVVVVVVVVREREREREREREVVVVREREREREREREVVVVREREVVVVVVVVREREVVVVZmZmREREREREVVVVVVVVREREREREVVVVREREVVVVVVVVZmZmVVVVVVVVVVVVREREREREREREREREREREREREVVVVREREVVVVVVVVVVVVVVVVREREREREREREREREREREVVVVREREVVVVREREREREREREVVVVREREREREREREVVVVREREREREMzMzREREVVVVREREREREMzMzREREREREZmZmd3d3mZmZu7u7qqqqiIiIREREMzMzMzMzVVVVVVVVMzMzMzMzIiIiMzMzMzMzREREVVVVREREIiIiMzMzREREVVVVMzMzIiIiERERIiIiERERERERIiIiERERIiIiIiIiMzMzIiIiIiIiIiIiMzMzIiIiVVVVVVVVREREMzMzREREVVVVREREMzMzMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREREREREREREREMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREMzMzREREREREREREREREREREMzMzREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzREREREREd3d3ZmZmREREREREREREREREREREMzMzMzMzMzMzREREMzMzREREVVVVREREZmZmVVVVVVVVd3d3ZmZmZmZmZmZmVVVVREREVVVVVVVVZmZmd3d3ZmZmVVVVVVVVVVVVVVVVZmZmd3d3ZmZmMzMzMzMzREREZmZmZmZmREREREREREREREREREREREREVVVVREREREREVVVVREREVVVVREREREREREREREREREREREREREREREREREREMzMzREREMzMzREREREREREREREREREREVVVVREREREREREREVVVVREREREREREREREREREREREREREREREREREREMzMzIiIiIiIiMzMzMzMzREREMzMzMzMzd3d3mZmZiIiIiIiId3d3ZmZmd3d3mZmZqqqqqqqqqqqqmZmZiIiIZmZmVVVVd3d3ZmZmZmZmZmZmZmZmVVVVZmZmZmZmd3d3iIiId3d3ZmZmd3d3qqqqu7u7mZmZiIiImZmZ3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////+7u7u7u7t3d3d3d3czMzN3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzN3d3czMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u8zMzLu7u7u7u6qqqru7u6qqqqqqqqqqqru7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqqqqqqqqqru7u6qqqru7u7u7u7u7u8zMzKqqqqqqqqqqqqqqqqqqqqqqqru7u7u7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqpmZmaqqqpmZmZmZmZmZmYiIiIiIiHd3d2ZmZmZmZlVVVVVVVURERERERERERERERERERDMzM0RERERERERERERERFVVVURERERERERERERERERERFVVVURERFVVVWZmZmZmZmZmZmZmZnd3d2ZmZnd3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZnd3d3d3d3d3d2ZmZmZmZnd3d3d3d2ZmZmZmZmZmZnd3d2ZmZlVVVWZmZlVVVWZmZnd3d2ZmZmZmZnd3d3d3d3d3d3d3d2ZmZlVVVURERDMzM1VVVWZmZkRERDMzM0RERERERERERERERERERFVVVVVVVURERFVVVURERERERCIiIjMzMzMzMzMzMzMzM0RERDMzM0RERFVVVURERERERERERFVVVURERERERERERFVVVURERERERDMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzM0RERERERERERDMzM0RERFVVVTMzM0RERDMzM0RERDMzMyIiIjMzMyIiIjMzMzMzMzMzMyIiIiIiIhERESIiIiIiIiIiIhERERERESIiIhERESIiIhERESIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzM0RERCIiIiIiIiIiIiIiIhERESIiIhERERERESIiIiIiIiIiIjMzM0RERERERFVVVWZmZkRERDMzMzMzM0RERDMzM0RERERERERERFVVVURERGZmZlVVVWZmZmZmZmZmZnd3d4iIiJmZmXd3d2ZmZlVVVVVVVURERGZmZlVVVURERFVVVVVVVURERERERERERERERDMzMzMzM0RERERERERERFVVVURERERERERERERERERERERERFVVVURERERERERERERERDMzM0RERDMzMzMzMzMzM0RERFVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZnd3d4iIiIiIiIiIiGZmZnd3d2ZmZlVVVWZmZnd3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZlVVVURERGZmZoiIiIiIiHd3d4iIiHd3d3d3d4iIiIiIiIiIiIiIiIiIiGZmZmZmZnd3d3d3d2ZmZkRERFVVVXd3d4iIiJmZmYiIiIiIiIiIiJmZmaqqqqqqqqqqqpmZmaqqqpmZmZmZmYiIiIiIiIiIiGZmZlVVVWZmZoiIiIiIiHd3d2ZmZoiIiHd3d3d3d3d3d5mZmYiIiIiIiHd3d2ZmZmZmZmZmZkRERFVVVVVVVURERFVVVVVVVVVVVXd3d5mZmYiIiHd3d4iIiHd3d4iIiIiIiIiIiIiIiHd3d2ZmZmZmZlVVVVVVVVVVVURERFVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVXd3d4iIiHd3d2ZmZmZmZnd3d2ZmZmZmZlVVVURERFVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d1VVVVVVVURERGZmZnd3d3d3d4iIiIiIiIiIiHd3d2ZmZlVVVVVVVURERERERERERERERERERERERERERERERFVVVURERERERDMzMzMzM0RERGZmZnd3d2ZmZlVVVURERFVVVURERFVVVVVVVVVVVURERERERERERERERERERERERFVVVVVVVVVVVTMzMzMzMzMzM1VVVXd3d4iIiHd3d1VVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVWZmZlVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVURERERERERERERERERERERERERERFVVVVVVVVVVVURERERERERERFVVVURERDMzM0RERGZmZlVVVVVVVVVVVWZmZmZmZlVVVVVVVURERERERDMzM0RERERERDMzM0RERDMzM0RERERERDMzM0RERERERDMzMzMzMzMzMzMzM0RERERERFVVVVVVVVVVVURERERERERERERERFVVVVVVVURERERERFVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVURERERERERERERERDMzMzMzMyIiIjMzMzMzM0RERERERDMzMzMzMzMzM0RERDMzM0RERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMyIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIhERERERESIiIiIiIiIiIiIiIkRERDMzMyIiIjMzM1VVVVVVVWZmZmZmZmZmZmZmZlVVVURERERERFVVVURERDMzM0RERERERERERERERERERERERFVVVURERERERFVVVWZmZlVVVVVVVVVVVURERERERERERERERERERERERFVVVWZmZmZmZmZmZlVVVURERDMzMzMzM0RERFVVVVVVVURERERERERERFVVVURERERERFVVVURERERERERERERERERERERERERERERERERERFVVVWZmZlVVVURERFVVVVVVVURERERERERERERERFVVVURERERERERERERERERERGZmZoiIiLu7u7u7u4iIiFVVVSIiIjMzMzMzM0RERDMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM0RERERERDMzMyIiIhERERERESIiIhERERERESIiIjMzM1VVVURERCIiIiIiIiIiIjMzMyIiIkRERFVVVURERDMzMzMzM1VVVURERDMzMyIiIiIiIjMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERDMzM0RERERERDMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERDMzM0RERDMzM0RERDMzM0RERDMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERDMzM0RERIiIiHd3d0RERERERERERERERDMzMzMzM0RERERERERERERERERERFVVVVVVVURERFVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVURERFVVVWZmZnd3d2ZmZlVVVWZmZmZmZmZmZnd3d3d3d1VVVSIiIkRERFVVVWZmZlVVVURERFVVVURERFVVVVVVVURERERERFVVVVVVVURERFVVVURERFVVVURERERERERERERERERERERERERERERERERERERERERERERERERERFVVVWZmZoiIiHd3d1VVVVVVVURERERERERERERERFVVVURERERERERERFVVVVVVVURERDMzMzMzMzMzMyIiIjMzMzMzM0RERDMzM1VVVZmZmZmZmYiIiIiIiHd3d3d3d5mZmaqqqpmZmaqqqru7u5mZmXd3d3d3d3d3d3d3d2ZmZnd3d2ZmZmZmZmZmZmZmZnd3d3d3d4iIiHd3d2ZmZoiIiLu7u7u7u6qqqpmZmaqqqt3d3e7u7v///+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////u7u7u7u7d3d3d3d3MzMzMzMzd3d3MzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3d3d3d3d3d3d3d3d3u7u7d3d3d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzd3d3MzMzMzMzd3d3MzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7vMzMy7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7uqqqq7u7u7u7u7u7vMzMy7u7u7u7u7u7u7u7u7u7uqqqqqqqqqqqq7u7u7u7u7u7u7u7uqqqqqqqqZmZmZmZmZmZmZmZmIiIiZmZmZmZmZmZmZmZmqqqqqqqqZmZmZmZmZmZmZmZmIiIh3d3d3d3dmZmZmZmZVVVVVVVVVVVVEREREREREREREREREREREREREREREREREREREREREREREREQzMzNERERERERERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3d3d3d3d3eIiIh3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3dmZmZ3d3d3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVmZmaIiIh3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3dmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVEREREREQzMzNERERVVVVVVVVVVVVmZmZVVVVmZmZVVVUzMzNEREREREREREQzMzMzMzNEREQzMzMiIiIzMzNVVVVVVVVVVVVEREQzMzNVVVVERERVVVVEREREREREREREREQzMzNEREQzMzMzMzNEREQzMzMzMzMiIiIzMzNVVVVVVVVEREREREREREQzMzNEREREREQzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzMzMzMiIiIiIiIREREiIiIiIiIiIiIiIiIiIiJEREQzMzMiIiIzMzMzMzMzMzNEREREREQiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMiIiIiIiIiIiIiIiIREREREREiIiIREREREREiIiIzMzMzMzMzMzNmZmaIiIhVVVVERERERERERERERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZ3d3eIiIh3d3dERERERERERERVVVVVVVVVVVVVVVVVVVVEREREREREREREREQzMzMzMzMzMzMzMzNERERERERVVVVVVVVVVVVERERERERVVVVERERVVVVEREREREQzMzNEREREREREREQzMzMzMzNVVVVVVVVmZmZ3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3eIiIiIiIh3d3dmZmZmZmZVVVVmZmZ3d3d3d3d3d3dmZmZmZmZmZmZ3d3eIiIh3d3d3d3d3d3dmZmZmZmZmZmZVVVVERERVVVWIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZmIiIiIiIiIiIiIiIhmZmZmZmZmZmZmZmZmZmZVVVVmZmaIiIiZmZmIiIiZmZmZmZmqqqqqqqqqqqqZmZmqqqqZmZmZmZmZmZmIiIiIiIiIiIhmZmZVVVV3d3d3d3eIiIh3d3d3d3d3d3eIiIh3d3d3d3eZmZmIiIh3d3d3d3d3d3dmZmZ3d3dVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZ3d3eZmZmIiIiIiIiIiIiIiIiZmZmZmZmIiIh3d3d3d3d3d3dmZmZERERERERERERERERVVVVVVVVmZmZmZmZmZmZmZmZERERVVVWIiIiIiIhmZmZ3d3d3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVERERVVVV3d3d3d3eZmZmZmZmIiIh3d3dmZmZmZmZmZmZVVVVVVVVEREQzMzNERERERERVVVVVVVVmZmZEREREREQzMzNERERVVVVVVVV3d3d3d3dmZmZVVVVERERVVVVERERVVVVVVVVVVVVERERERERERERERERERERVVVVVVVVEREQzMzMzMzMzMzNVVVV3d3d3d3eIiIhmZmZVVVVVVVVVVVVmZmZVVVVmZmZVVVVmZmZVVVVmZmZmZmZmZmZmZmZVVVVVVVVERERERERERERVVVVVVVVmZmZVVVVVVVVVVVVERERERERVVVVVVVVVVVVERERVVVVVVVVVVVVERERERERVVVVERERERERERERmZmZmZmZmZmZVVVVVVVVmZmZmZmZEREREREREREREREQzMzMzMzNEREREREQzMzNEREREREREREREREREREQzMzNEREQzMzMzMzNERERVVVVERERVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVERERERERVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVERERERERVVVVEREQzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMiIiIiIiIzMzMiIiIiIiIiIiIiIiIREREiIiIREREREREiIiIiIiIREREiIiIiIiIiIiIzMzMiIiIzMzNVVVVVVVVmZmZmZmZmZmZVVVVERERVVVVEREREREREREQzMzMzMzNEREREREREREREREREREREREREREQzMzNERERVVVVVVVVERERVVVVVVVVEREREREQzMzNEREQzMzNVVVVVVVVVVVVERERERERERERERERERERERERVVVVVVVVERERERERERERERERVVVVEREREREREREREREREREREREREREQzMzMzMzNERERVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERVVVVERERVVVVVVVV3d3eZmZl3d3dEREQiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIzMzNEREREREREREQzMzNEREREREREREQzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzNEREREREQiIiIzMzMiIiIzMzMzMzMiIiJERERERERERERERERmZmZEREREREQiIiIzMzMiIiIzMzMzMzMzMzMzMzNEREQzMzNEREREREQzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNEREREREREREREREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzMiIiIzMzMiIiIzMzMzMzNVVVVEREREREQzMzNERER3d3eZmZlVVVVERERERERERERERERERERERERVVVVERERERERERERERERVVVVVVVVERERERERmZmZmZmZmZmZmZmZVVVVERERVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVmZmZ3d3dmZmYzMzMzMzNVVVV3d3dmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVERERERERERERERERERERVVVV3d3dVVVVERERERERERERVVVVVVVVVVVVVVVVmZmaIiIh3d3dVVVVVVVVERERVVVVERERVVVVERERERERVVVVERERVVVVVVVVVVVUzMzMzMzMzMzMzMzMzMzNEREQzMzNEREQzMzN3d3eZmZmIiIiIiIiZmZl3d3eZmZmqqqqqqqqqqqqqqqqZmZmIiIh3d3d3d3dmZmZVVVVVVVVmZmZmZmZmZmZVVVV3d3dmZmZ3d3eIiIh3d3dmZmaIiIi7u7u7u7uqqqqZmZmqqqrMzMzu7u7u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////7u7u7u7uzMzMu7u7u7u7u7u7u7u7u7u7u7u7zMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM3d3d3d3d3d3dzMzM3d3d3d3d3d3d3d3dzMzM3d3d3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7zMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7zMzMu7u7u7u7zMzMu7u7u7u7u7u7qqqqu7u7u7u7u7u7qqqqu7u7qqqqu7u7qqqqqqqqqqqqqqqqmZmZmZmZmZmZmZmZmZmZmZmZiIiImZmZmZmZqqqqmZmZmZmZmZmZmZmZmZmZiIiIiIiIiIiId3d3d3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVREREREREREREVVVVVVVVREREVVVVVVVVREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3d3d3iIiId3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3iIiId3d3d3d3iIiIiIiImZmZiIiId3d3iIiId3d3ZmZmVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmVVVVZmZmd3d3d3d3ZmZmVVVVVVVVREREREREVVVVREREREREZmZmZmZmZmZmZmZmVVVVREREMzMzMzMzREREREREVVVVREREREREMzMzMzMzVVVVZmZmREREREREMzMzREREVVVVVVVVVVVVREREREREMzMzIiIiMzMzMzMzMzMzREREREREMzMzMzMzMzMzVVVVZmZmVVVVVVVVREREREREMzMzMzMzMzMzMzMzVVVVREREREREMzMzMzMzMzMzMzMzMzMzREREREREMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiERERIiIiREREMzMzMzMzREREZmZmREREMzMzIiIiIiIiMzMzMzMzREREREREREREREREREREMzMzVVVVVVVVVVVVVVVVVVVVMzMzIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiMzMzMzMzZmZmiIiIZmZmREREMzMzREREVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3d3d3d3d3VVVVVVVVVVVVVVVVVVVVZmZmVVVVREREREREREREREREREREVVVVVVVVVVVVREREREREREREREREREREMzMzIiIiMzMzREREd3d3VVVVREREVVVVVVVVVVVVVVVVREREVVVVREREREREREREVVVVREREREREREREREREVVVVd3d3iIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiId3d3ZmZmVVVVZmZmZmZmd3d3d3d3d3d3ZmZmd3d3ZmZmd3d3d3d3d3d3d3d3ZmZmd3d3VVVVVVVVREREREREd3d3mZmZiIiIiIiImZmZmZmZiIiIiIiIiIiIiIiId3d3iIiId3d3ZmZmZmZmZmZmZmZmZmZmd3d3d3d3iIiImZmZmZmZqqqqqqqqmZmZiIiImZmZqqqqmZmZmZmZmZmZiIiId3d3VVVVVVVVZmZmd3d3d3d3d3d3iIiImZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3ZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmmZmZmZmZmZmZmZmZmZmZiIiImZmZiIiId3d3d3d3ZmZmVVVVREREREREVVVVVVVVVVVVVVVVZmZmd3d3ZmZmZmZmREREVVVVZmZmiIiIiIiId3d3d3d3d3d3ZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmd3d3ZmZmZmZmVVVVZmZmiIiIiIiIiIiImZmZd3d3d3d3ZmZmVVVVVVVVZmZmVVVVMzMzREREREREVVVVVVVVVVVVVVVVVVVVREREMzMzREREVVVVZmZmd3d3d3d3ZmZmVVVVREREREREVVVVVVVVVVVVVVVVVVVVREREREREVVVVREREVVVVVVVVREREREREREREMzMzREREZmZmd3d3iIiId3d3ZmZmVVVVZmZmZmZmVVVVVVVVZmZmVVVVZmZmZmZmd3d3ZmZmZmZmVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREVVVVREREREREVVVVVVVVVVVVREREVVVVREREREREREREREREVVVVZmZmd3d3VVVVVVVVZmZmVVVVREREREREREREMzMzREREREREMzMzREREREREREREREREREREVVVVVVVVREREREREMzMzMzMzVVVVVVVVREREVVVVVVVVREREVVVVREREREREVVVVREREREREVVVVVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVREREREREREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREREREVVVVVVVVREREREREREREMzMzREREREREMzMzMzMzMzMzMzMzREREREREREREMzMzIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERERERIiIiIiIiIiIiIiIiIiIiMzMzREREVVVVZmZmZmZmZmZmVVVVVVVVREREREREREREMzMzREREREREMzMzREREREREREREREREREREMzMzREREMzMzMzMzREREVVVVREREREREREREREREREREMzMzREREREREREREVVVVREREREREREREMzMzREREREREREREMzMzMzMzREREREREVVVVVVVVZmZmVVVVREREREREMzMzREREMzMzMzMzMzMzREREREREREREVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREVVVVVVVVREREREREREREREREVVVVREREREREMzMzIiIiERERIiIiERERIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzIiIiMzMzMzMzIiIiMzMzIiIiMzMzMzMzREREVVVVVVVVVVVVMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREREREREREREREREREREREREREVVVVVVVVREREREREMzMzMzMzMzMzMzMzREREMzMzMzMzIiIiMzMzMzMzMzMzMzMzREREZmZmVVVVREREMzMzMzMzZmZmd3d3REREREREMzMzREREREREREREREREREREREREREREREREREREZmZmZmZmVVVVVVVVZmZmd3d3ZmZmd3d3VVVVREREREREVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVZmZmVVVVIiIiREREZmZmiIiIZmZmVVVVREREVVVVVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREVVVVZmZmiIiIZmZmREREREREREREREREREREREREREREREREVVVVVVVVREREVVVVVVVVREREVVVVZmZmZmZmVVVVREREVVVVVVVVVVVVREREREREMzMzMzMzMzMzREREREREREREREREMzMzVVVVmZmZqqqqmZmZmZmZiIiIiIiImZmZmZmZmZmZiIiId3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmiIiImZmZu7u7u7u7mZmZqqqq3d3d7u7u7u7u7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////+7u7t3d3bu7u7u7u7u7u8zMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzN3d3czMzMzMzN3d3czMzN3d3czMzMzMzMzMzMzMzN3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3czMzMzMzMzMzLu7u7u7u8zMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u8zMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u8zMzLu7u7u7u7u7u8zMzLu7u7u7u8zMzMzMzLu7u8zMzLu7u6qqqru7u7u7u7u7u7u7u7u7u7u7u6qqqru7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqpmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiJmZmZmZmZmZmaqqqpmZmZmZmYiIiJmZmYiIiIiIiHd3d3d3d2ZmZlVVVWZmZlVVVURERFVVVURERFVVVVVVVURERFVVVVVVVVVVVURERFVVVVVVVURERERERERERERERERERERERFVVVVVVVWZmZlVVVWZmZmZmZnd3d4iIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiHd3d4iIiJmZmYiIiIiIiHd3d3d3d4iIiHd3d2ZmZmZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d2ZmZmZmZlVVVWZmZmZmZlVVVVVVVVVVVURERFVVVWZmZoiIiHd3d1VVVURERERERFVVVVVVVVVVVURERERERERERGZmZlVVVURERERERERERDMzM0RERHd3d2ZmZlVVVURERDMzMyIiIjMzMzMzMzMzM0RERERERDMzMzMzMyIiIkRERFVVVWZmZlVVVVVVVURERERERERERERERERERFVVVWZmZlVVVURERERERERERDMzMzMzM1VVVVVVVTMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMyIiIiIiIjMzM1VVVURERERERERERFVVVTMzMzMzMzMzMzMzM0RERERERERERFVVVVVVVVVVVURERERERFVVVWZmZmZmZlVVVURERERERDMzMzMzM0RERERERDMzMyIiIjMzMyIiIiIiIhERESIiIiIiIiIiIhERESIiIjMzM0RERFVVVWZmZlVVVVVVVURERFVVVVVVVVVVVWZmZnd3d2ZmZmZmZmZmZnd3d3d3d2ZmZmZmZlVVVURERERERERERGZmZmZmZlVVVVVVVURERFVVVVVVVVVVVWZmZlVVVVVVVURERFVVVURERERERERERDMzMzMzM0RERHd3d3d3d1VVVVVVVVVVVWZmZkRERFVVVVVVVURERFVVVVVVVVVVVURERERERERERERERGZmZmZmZnd3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d2ZmZlVVVWZmZnd3d2ZmZmZmZnd3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZlVVVURERERERHd3d5mZmZmZmYiIiJmZmZmZmYiIiIiIiIiIiJmZmYiIiIiIiIiIiHd3d3d3d1VVVWZmZmZmZmZmZnd3d5mZmZmZmZmZmZmZmZmZmYiIiJmZmZmZmaqqqpmZmZmZmYiIiHd3d2ZmZmZmZmZmZmZmZmZmZnd3d3d3d5mZmZmZmXd3d4iIiJmZmYiIiIiIiIiIiIiIiIiIiGZmZmZmZmZmZlVVVWZmZmZmZnd3d1VVVVVVVVVVVWZmZmZmZmZmZpmZmZmZmaqqqpmZmYiIiIiIiIiIiHd3d2ZmZmZmZlVVVVVVVVVVVVVVVURERFVVVVVVVWZmZnd3d2ZmZlVVVURERERERFVVVXd3d4iIiJmZmXd3d2ZmZlVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVWZmZmZmZnd3d3d3d1VVVVVVVWZmZoiIiJmZmYiIiIiIiHd3d2ZmZmZmZlVVVWZmZmZmZlVVVURERFVVVVVVVVVVVURERGZmZlVVVURERERERDMzMzMzM0RERGZmZnd3d3d3d2ZmZlVVVVVVVURERERERERERFVVVWZmZlVVVURERFVVVVVVVVVVVVVVVURERERERERERDMzM0RERFVVVWZmZnd3d2ZmZnd3d2ZmZmZmZmZmZlVVVWZmZlVVVWZmZmZmZmZmZnd3d3d3d3d3d2ZmZlVVVVVVVVVVVURERERERFVVVVVVVVVVVWZmZlVVVVVVVVVVVURERERERFVVVURERFVVVURERFVVVURERFVVVURERFVVVURERERERDMzMzMzM1VVVWZmZmZmZlVVVVVVVVVVVURERERERERERDMzMzMzMzMzM0RERERERDMzM0RERFVVVURERFVVVVVVVVVVVURERDMzMzMzM1VVVVVVVURERERERFVVVVVVVURERFVVVURERFVVVURERERERERERFVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERDMzMyIiIjMzMzMzMzMzM0RERERERERERDMzM0RERERERDMzM0RERDMzM0RERERERDMzMyIiIiIiIjMzMyIiIjMzM0RERERERCIiIjMzMyIiIiIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIjMzMzMzM0RERFVVVURERFVVVVVVVWZmZlVVVURERDMzMzMzM0RERERERERERERERERERERERERERERERERERDMzM0RERDMzM0RERERERFVVVURERERERERERERERDMzM0RERERERERERERERERERERERDMzM0RERDMzM0RERERERERERERERERERFVVVVVVVVVVVWZmZlVVVVVVVTMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERFVVVWZmZmZmZlVVVURERERERERERFVVVWZmZlVVVURERDMzM0RERERERERERDMzMzMzMyIiIiIiIiIiIhERESIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzM0RERDMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERDMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVURERDMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzM0RERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERFVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVURERERERDMzMzMzM0RERGZmZlVVVURERERERERERERERERERERERERERDMzMzMzM0RERERERFVVVVVVVURERFVVVWZmZnd3d2ZmZmZmZlVVVURERFVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVWZmZmZmZkRERDMzM0RERGZmZmZmZmZmZlVVVWZmZlVVVWZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZlVVVWZmZlVVVURERERERFVVVWZmZnd3d2ZmZkRERDMzM0RERDMzM0RERDMzM0RERERERDMzM0RERERERFVVVURERERERFVVVVVVVXd3d2ZmZlVVVVVVVVVVVURERERERERERERERERERDMzMzMzM0RERERERERERERERERERERERHd3d6qqqpmZmYiIiIiIiHd3d4iIiJmZmXd3d3d3d3d3d2ZmZmZmZlVVVURERGZmZmZmZkRERFVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d4iIiIiIiKqqqqqqqru7u8zMzN3d3d3d3d3d3e7u7v///////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3u7u7u7u7d3d3u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3MzMzd3d3MzMzMzMzMzMzMzMy7u7vMzMzMzMzMzMy7u7u7u7uqqqq7u7uqqqqqqqq7u7uqqqq7u7u7u7vMzMy7u7vMzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7uqqqq7u7u7u7u7u7u7u7u7u7u7u7u7u7uqqqq7u7uqqqqqqqqqqqqqqqqqqqqZmZmqqqqZmZmZmZmZmZmIiIiZmZmZmZmZmZmIiIiZmZmZmZmIiIiZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmIiIiIiIh3d3dmZmZmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVERERVVVVVVVVmZmZmZmZmZmZmZmZ3d3d3d3dmZmZ3d3eIiIh3d3eIiIh3d3eIiIh3d3d3d3d3d3eIiIiZmZmIiIiIiIiIiIiIiIiIiIh3d3eIiIiIiIiIiIiIiIh3d3dVVVVVVVVmZmZ3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZ3d3d3d3dVVVVmZmZVVVVmZmZ3d3eIiIhmZmZVVVVERERERER3d3dmZmZVVVVVVVVVVVVVVVVmZmZEREQzMzNEREREREREREQzMzN3d3eIiIhVVVUzMzNEREQzMzMzMzMzMzNEREQzMzMzMzNEREREREQzMzNERERVVVVVVVUzMzNVVVVVVVVmZmZVVVVERERVVVVmZmZmZmZ3d3dmZmZVVVVERERERERVVVVmZmZEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERVVVVVVVVVVVVEREQzMzMzMzNERERERERERERERERmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVEREQzMzNEREREREREREQzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIREREREREiIiIzMzNERERVVVVmZmZmZmZ3d3dmZmZVVVVVVVVmZmZmZmZ3d3dmZmZmZmZmZmZ3d3d3d3dmZmZmZmZmZmZERERVVVVVVVVmZmZmZmZVVVVERERVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVERERERERERERERERERERVVVVVVVVmZmaIiIhmZmZVVVVmZmZmZmZVVVVVVVVVVVVmZmZVVVVVVVVmZmZVVVVEREQzMzNERERVVVVmZmZmZmZmZmZ3d3d3d3d3d3eZmZmZmZmZmZmZmZmqqqqZmZmIiIiIiIhVVVVmZmZ3d3d3d3d3d3dmZmZVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZERERERERVVVWZmZmZmZmZmZmIiIiZmZmIiIiIiIiZmZmIiIiZmZl3d3eIiIiIiIhVVVVVVVVmZmZ3d3dmZmZ3d3eZmZmZmZmIiIiIiIiZmZmZmZmqqqqZmZmqqqqZmZmIiIh3d3dmZmZ3d3dmZmZ3d3dmZmZmZmZ3d3eIiIiZmZmZmZmIiIiZmZmIiIiIiIiIiIiZmZl3d3eIiIh3d3d3d3d3d3dVVVVmZmZ3d3d3d3dmZmZmZmZmZmZmZmZVVVVmZmZmZmaIiIiZmZmZmZl3d3eIiIiZmZmIiIhmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVV3d3d3d3dVVVVEREQzMzNERERmZmaIiIiZmZl3d3dVVVVVVVVERERVVVVmZmZmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZVVVV3d3eZmZmIiIiIiIh3d3dmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVEREREREQzMzMzMzNERER3d3eIiIh3d3dVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVEREREREREREREREQzMzNERERmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dVVVVVVVVVVVVERERERERERERVVVVmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVERERVVVVERERERERVVVVVVVVERERERERVVVVEREREREQzMzNERERVVVVmZmZmZmZVVVVVVVVmZmZVVVVERERVVVVEREREREREREREREREREQzMzNERERERERERERERERVVVVEREREREREREQzMzNERERVVVVERERVVVVERERERERERERVVVVVVVVVVVVERERERERERERVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVERERVVVVERERERERVVVVmZmZVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREREREREREQzMzMzMzNEREQzMzNEREQzMzMzMzMiIiIiIiIzMzMiIiJEREQzMzMzMzMzMzMiIiIREREiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzNERERVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERVVVVVVVVERERERERERERVVVVVVVVEREREREQzMzNEREREREQzMzNEREREREREREREREQzMzNEREQzMzNEREREREREREREREQzMzNEREQzMzNEREQzMzMzMzMzMzNVVVVmZmZmZmZVVVVVVVVVVVVEREQzMzNEREQzMzNERERERERERERERERERERERERERERVVVVVVVVVVVVERERERERERERERERERERVVVUzMzMzMzNEREREREQzMzMiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMiIiIzMzNEREREREQzMzMzMzNEREQzMzNEREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzNERERVVVVEREREREQzMzMzMzNEREQzMzNEREQzMzNEREQzMzNERERERERERERVVVVERERVVVVVVVVVVVVERERVVVVVVVVERERERERERERVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVVVVVVVVUzMzMzMzNERERERERVVVVmZmZERERVVVVEREREREREREQzMzNEREQzMzMzMzMzMzNERERERERERERVVVVVVVVmZmZ3d3d3d3dVVVVVVVVERERVVVVVVVVmZmZmZmZmZmZVVVVmZmZmZmZ3d3dmZmYzMzMzMzNmZmaIiIh3d3dmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZVVVVmZmZmZmZ3d3d3d3d3d3dmZmZmZmZmZmZVVVVmZmZVVVUzMzMzMzNEREQzMzNEREREREREREREREQzMzNEREREREQzMzNERERERERERERERERVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVEREREREQzMzNERER3d3eIiIhEREREREQzMzNmZmaZmZmqqqqZmZmZmZmIiIh3d3eIiIiIiIh3d3d3d3d3d3d3d3dVVVVVVVVmZmZVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3d3d3eIiIiqqqq7u7vMzMzMzMzd3d3d3d3d3d3u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////7u7u////////////////////7u7u7u7u3d3d7u7u7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u3d3d7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7zMzMzMzMzMzMzMzMzMzM3d3dzMzMzMzMzMzMzMzMzMzMu7u7u7u7zMzMu7u7u7u7u7u7zMzMzMzMu7u7u7u7u7u7qqqqqqqqqqqqu7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqmZmZmZmZmZmZmZmZiIiImZmZmZmZmZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZmZmZmZmZmZmZiIiIiIiImZmZiIiIiIiIiIiIiIiIZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVZmZmVVVVREREREREVVVVZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmd3d3d3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3mZmZiIiIiIiId3d3ZmZmVVVVZmZmd3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmiIiId3d3d3d3d3d3ZmZmd3d3ZmZmd3d3ZmZmZmZmVVVVVVVVVVVVd3d3ZmZmiIiId3d3ZmZmVVVVZmZmZmZmREREVVVVVVVVREREREREVVVViIiId3d3VVVVREREREREVVVVVVVVREREREREMzMzMzMzVVVVREREREREVVVVVVVVREREREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmREREZmZmd3d3ZmZmZmZmREREVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzVVVVREREZmZmZmZmVVVVZmZmREREREREVVVVVVVVZmZmVVVVZmZmd3d3d3d3VVVVd3d3ZmZmVVVVVVVVREREVVVVREREMzMzREREVVVVREREMzMzIiIiIiIiIiIiIiIiIiIiREREREREIiIiIiIiMzMzREREVVVVVVVVZmZmZmZmd3d3d3d3ZmZmZmZmVVVVZmZmd3d3ZmZmd3d3d3d3d3d3d3d3iIiIZmZmZmZmVVVVREREREREVVVVZmZmZmZmVVVVZmZmVVVVVVVVZmZmZmZmVVVVREREVVVVVVVVVVVVVVVVREREREREREREVVVVZmZmd3d3ZmZmZmZmZmZmZmZmd3d3ZmZmZmZmVVVVVVVVREREVVVVVVVVVVVVREREREREREREZmZmd3d3d3d3d3d3d3d3d3d3iIiIqqqqmZmZiIiIqqqqqqqqiIiId3d3ZmZmZmZmd3d3d3d3ZmZmZmZmZmZmd3d3iIiIiIiIiIiIiIiIiIiIiIiIZmZmVVVVd3d3iIiIVVVVREREVVVViIiImZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmVVVVVVVVZmZmZmZmd3d3ZmZmd3d3mZmZqqqqqqqqmZmZqqqqmZmZqqqqmZmZiIiIiIiId3d3d3d3ZmZmZmZmZmZmd3d3d3d3d3d3d3d3iIiIqqqqqqqqmZmZmZmZmZmZiIiIiIiIiIiImZmZiIiId3d3ZmZmVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmd3d3iIiImZmZmZmZiIiId3d3ZmZmVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVZmZmd3d3d3d3ZmZmREREREREVVVVd3d3iIiImZmZd3d3ZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3ZmZmVVVVZmZmiIiIiIiIiIiId3d3d3d3ZmZmZmZmVVVVREREREREZmZmVVVVZmZmVVVVVVVVZmZmVVVVVVVVREREMzMzMzMzZmZmd3d3iIiIiIiIZmZmVVVVVVVVREREREREREREVVVVREREVVVVREREVVVVVVVVVVVVREREREREREREMzMzREREMzMzZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3ZmZmVVVVVVVVREREVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVREREREREVVVVREREVVVVREREVVVVVVVVREREREREVVVVZmZmZmZmZmZmVVVVZmZmVVVVREREVVVVREREREREREREREREREREREREREREREREVVVVREREREREVVVVREREREREREREREREVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVREREREREVVVVVVVVREREVVVVVVVVVVVVVVVVREREVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmVVVVMzMzREREREREREREMzMzMzMzREREMzMzREREREREREREREREREREMzMzMzMzREREREREREREREREREREMzMzMzMzMzMzIiIiIiIiERERMzMzREREMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiIiIiVVVVVVVVVVVVZmZmVVVVREREREREREREVVVVVVVVZmZmVVVVVVVVVVVVREREREREREREREREREREREREREREREREMzMzMzMzVVVVVVVVREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREZmZmVVVVREREREREMzMzREREMzMzVVVVREREREREREREREREREREREREREREREREVVVVVVVVREREVVVVREREREREREREREREVVVVREREMzMzMzMzMzMzIiIiIiIiMzMzIiIiERERIiIiIiIiMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREMzMzMzMzMzMzVVVVVVVVREREREREREREMzMzMzMzREREVVVVVVVVMzMzIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzREREREREVVVVVVVVREREREREVVVVREREREREREREREREREREREREREREVVVVREREREREVVVVREREVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzVVVVVVVVREREREREMzMzREREREREREREVVVVVVVVREREVVVVREREREREREREMzMzREREMzMzREREMzMzREREREREREREVVVVZmZmd3d3iIiId3d3REREREREVVVVREREZmZmVVVVZmZmZmZmVVVVZmZmd3d3VVVVIiIiREREiIiImZmZiIiId3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmZmZmd3d3ZmZmd3d3d3d3ZmZmREREREREMzMzREREREREREREMzMzREREREREREREVVVVVVVVREREREREVVVVREREVVVVREREREREVVVVREREVVVVVVVVVVVVVVVVZmZmVVVVREREREREREREREREREREREREd3d3qqqqd3d3VVVVREREREREd3d3qqqqmZmZmZmZmZmZmZmZmZmZd3d3d3d3d3d3qqqqmZmZd3d3ZmZmZmZmZmZmVVVVREREVVVVREREVVVVREREREREREREVVVVVVVVZmZmZmZmZmZmZmZmd3d3iIiImZmZqqqqu7u7u7u7zMzM3d3d3d3d3d3d7u7u7u7u////////////7u7u////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////+7u7u7u7u7u7t3d3czMzMzMzMzMzMzMzN3d3czMzLu7u7u7u7u7u7u7u7u7u8zMzN3d3czMzN3d3czMzMzMzLu7u7u7u8zMzLu7u7u7u7u7u6qqqru7u6qqqru7u6qqqru7u7u7u7u7u7u7u8zMzMzMzMzMzMzMzMzMzMzMzLu7u8zMzMzMzLu7u8zMzLu7u7u7u8zMzLu7u8zMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u8zMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u8zMzLu7u8zMzLu7u6qqqru7u6qqqqqqqqqqqqqqqqqqqpmZmZmZmYiIiJmZmZmZmaqqqpmZmZmZmZmZmYiIiJmZmYiIiJmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiHd3d3d3d3d3d4iIiHd3d4iIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiJmZmYiIiIiIiJmZmYiIiIiIiIiIiIiIiHd3d3d3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVWZmZnd3d2ZmZlVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d2ZmZmZmZoiIiIiIiGZmZmZmZnd3d3d3d3d3d4iIiHd3d2ZmZnd3d4iIiHd3d2ZmZnd3d4iIiHd3d3d3d3d3d3d3d2ZmZmZmZlVVVVVVVWZmZmZmZpmZmZmZmXd3d1VVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVYiIiIiIiFVVVURERFVVVVVVVWZmZlVVVURERERERDMzM0RERFVVVWZmZnd3d3d3d3d3d1VVVURERERERGZmZnd3d3d3d3d3d2ZmZlVVVVVVVURERFVVVXd3d3d3d3d3d3d3d2ZmZmZmZlVVVURERERERERERERERERERERERERERFVVVVVVVURERFVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVWZmZmZmZkRERERERERERFVVVURERERERDMzMzMzMyIiIiIiIjMzM1VVVURERDMzMyIiIjMzM0RERFVVVVVVVWZmZnd3d3d3d3d3d3d3d3d3d1VVVWZmZnd3d3d3d4iIiHd3d4iIiIiIiHd3d2ZmZlVVVVVVVVVVVVVVVVVVVXd3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZlVVVURERFVVVVVVVXd3d3d3d2ZmZnd3d3d3d4iIiHd3d2ZmZmZmZlVVVVVVVVVVVURERFVVVVVVVVVVVTMzM1VVVWZmZnd3d4iIiIiIiIiIiIiIiIiIiJmZmZmZmYiIiJmZmYiIiIiIiIiIiGZmZmZmZmZmZnd3d4iIiIiIiHd3d4iIiIiIiJmZmZmZmYiIiHd3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d2ZmZlVVVXd3d5mZmZmZmZmZmYiIiIiIiIiIiIiIiHd3d3d3d2ZmZlVVVWZmZnd3d2ZmZnd3d3d3d3d3d4iIiKqqqru7u7u7u6qqqqqqqqqqqpmZmYiIiIiIiIiIiHd3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d3d3d4iIiKqqqqqqqqqqqqqqqoiIiJmZmXd3d3d3d4iIiIiIiHd3d2ZmZlVVVWZmZnd3d2ZmZmZmZmZmZmZmZnd3d3d3d2ZmZlVVVVVVVXd3d5mZmaqqqqqqqpmZmXd3d2ZmZlVVVURERFVVVWZmZnd3d1VVVVVVVVVVVWZmZnd3d3d3d2ZmZlVVVURERGZmZnd3d5mZmYiIiHd3d3d3d3d3d2ZmZnd3d3d3d4iIiHd3d3d3d4iIiIiIiHd3d3d3d3d3d2ZmZnd3d1VVVWZmZoiIiIiIiIiIiIiIiHd3d2ZmZlVVVVVVVURERERERFVVVVVVVWZmZnd3d2ZmZlVVVVVVVVVVVURERDMzM0RERGZmZoiIiIiIiIiIiGZmZlVVVVVVVURERFVVVVVVVVVVVVVVVURERFVVVVVVVVVVVURERERERERERDMzMzMzM0RERERERFVVVWZmZmZmZmZmZmZmZlVVVVVVVWZmZnd3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZlVVVURERFVVVVVVVVVVVWZmZnd3d2ZmZlVVVVVVVVVVVVVVVURERERERERERFVVVVVVVURERERERERERERERFVVVURERERERERERFVVVVVVVXd3d2ZmZmZmZmZmZlVVVVVVVURERFVVVURERERERERERFVVVURERERERERERFVVVURERERERFVVVVVVVURERERERDMzM2ZmZmZmZlVVVVVVVVVVVVVVVVVVVURERFVVVURERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVURERFVVVVVVVXd3d1VVVURERERERFVVVURERDMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERDMzMzMzM0RERERERERERERERERERCIiIjMzMyIiIiIiIiIiIjMzM0RERDMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzM1VVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVURERDMzMzMzMzMzMzMzM0RERERERERERERERFVVVVVVVVVVVURERERERDMzM0RERDMzM0RERERERDMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM1VVVVVVVURERDMzM0RERERERERERERERERERERERERERERERERERDMzM0RERFVVVWZmZlVVVURERERERERERFVVVVVVVURERFVVVVVVVTMzMyIiIjMzMyIiIjMzMzMzMyIiIiIiIiIiIkRERERERERERERERERERDMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERERERERERDMzMzMzMyIiIkRERERERERERDMzMzMzMzMzM0RERERERFVVVVVVVURERDMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERERERERERERERERERERERFVVVVVVVVVVVURERERERERERFVVVURERFVVVURERERERERERERERERERERERERERERERFVVVVVVVVVVVVVVVURERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERGZmZkRERERERERERERERDMzM0RERFVVVVVVVURERERERERERERERERERDMzM0RERDMzMzMzM0RERERERERERFVVVURERFVVVXd3d3d3d1VVVURERFVVVURERFVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d1VVVTMzM2ZmZqqqqru7u7u7u5mZmXd3d3d3d3d3d2ZmZnd3d2ZmZmZmZmZmZlVVVWZmZmZmZlVVVVVVVWZmZmZmZlVVVURERERERFVVVURERERERERERFVVVVVVVWZmZmZmZnd3d1VVVVVVVVVVVURERFVVVVVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVWZmZnd3d1VVVVVVVURERERERERERERERFVVVZmZmZmZmWZmZlVVVTMzM2ZmZqqqqqqqqqqqqqqqqpmZmYiIiHd3d1VVVWZmZqqqqru7u6qqqnd3d3d3d5mZmXd3d2ZmZlVVVURERERERFVVVURERERERFVVVURERFVVVVVVVWZmZmZmZnd3d4iIiIiIiKqqqqqqqru7u7u7u8zMzN3d3bu7u8zMzO7u7v///////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////u7u7////////////////////////////////MzMzMzMy7u7u7u7u7u7uqqqq7u7uqqqq7u7u7u7u7u7uqqqqZmZmZmZmqqqqqqqqqqqqqqqqZmZmqqqqqqqqqqqqqqqqqqqqZmZmZmZmIiIiIiIiIiIh3d3d3d3d3d3d3d3eIiIiIiIiIiIiZmZmZmZmZmZmZmZmqqqqZmZmqqqqqqqq7u7uqqqqZmZmZmZmZmZmZmZmqqqqZmZmZmZmZmZmqqqqqqqqqqqq7u7uqqqq7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7vMzMy7u7u7u7u7u7u7u7u7u7vMzMy7u7u7u7u7u7vMzMy7u7uqqqq7u7u7u7uqqqqqqqqqqqqqqqqZmZmqqqqZmZmqqqqIiIiZmZmZmZmZmZmZmZmZmZmZmZmqqqqqqqqZmZmZmZmZmZmIiIiIiIiIiIiIiIh3d3d3d3eIiIh3d3d3d3d3d3d3d3eIiIh3d3eIiIh3d3eIiIiIiIh3d3eIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIh3d3eIiIiIiIhmZmZmZmZmZmZmZmZVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVmZmZ3d3d3d3dmZmZmZmZVVVVVVVVmZmZVVVVERERERERVVVVERERERERVVVVERERVVVVmZmZ3d3d3d3d3d3dmZmZ3d3d3d3dmZmZmZmZmZmZ3d3d3d3d3d3eIiIiIiIh3d3dmZmZmZmZ3d3d3d3eIiIh3d3dVVVV3d3eZmZl3d3dVVVV3d3eIiIh3d3d3d3d3d3d3d3d3d3dmZmZVVVVVVVVmZmZmZmaIiIiZmZlmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZ3d3eIiIhmZmZVVVVVVVVVVVVmZmZVVVVVVVVERERERERERERVVVWIiIiIiIiIiIh3d3dmZmZVVVVVVVV3d3d3d3d3d3d3d3dmZmZmZmZVVVVmZmZVVVV3d3d3d3dmZmZmZmZ3d3d3d3d3d3dVVVVVVVVmZmZmZmZVVVVVVVVVVVVmZmZmZmZVVVVERERmZmZmZmZ3d3dmZmaIiIhmZmZmZmZmZmZ3d3d3d3d3d3d3d3eIiIh3d3dmZmZmZmZ3d3dmZmZmZmZVVVUzMzNERERVVVVVVVVEREREREQiIiIzMzMiIiJERERmZmZEREQzMzMzMzMzMzNERERERERVVVVmZmZ3d3d3d3d3d3d3d3eIiIiIiIh3d3dmZmZmZmaIiIiZmZmIiIiZmZmIiIhmZmZVVVVmZmZVVVVVVVV3d3dmZmZVVVVmZmZ3d3dmZmZmZmZVVVVVVVVmZmZ3d3d3d3d3d3dmZmZmZmZVVVVERERERERVVVVmZmZmZmZ3d3d3d3eIiIiIiIiIiIhmZmZmZmZVVVVERERERERVVVVVVVVVVVVVVVVERERVVVVmZmaIiIiIiIiIiIiIiIiZmZmZmZmZmZmIiIiIiIiZmZl3d3eIiIiIiIhmZmZmZmZmZmZ3d3eIiIiIiIiIiIh3d3d3d3eIiIiIiIiIiIiIiIiIiIhmZmZmZmZVVVVVVVVmZmZmZmZmZmZVVVV3d3eZmZmZmZmqqqqqqqqZmZmZmZmIiIiIiIh3d3d3d3dmZmZ3d3d3d3d3d3dmZmZ3d3eIiIiIiIiIiIiqqqq7u7u7u7u7u7uqqqqZmZmZmZmIiIh3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3dmZmZ3d3eZmZmqqqqZmZmqqqqqqqqZmZmIiIh3d3d3d3eIiIh3d3d3d3dmZmZVVVV3d3d3d3dmZmZ3d3d3d3dmZmZ3d3eIiIhmZmZVVVVVVVVVVVV3d3eZmZmZmZmIiIh3d3dmZmZmZmZVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZ3d3eIiIh3d3dVVVVVVVVmZmaIiIiIiIiIiIiIiIh3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIh3d3dmZmZmZmZ3d3d3d3eIiIiZmZmIiIiIiIh3d3dmZmZVVVVERERVVVVERERVVVVmZmZmZmZ3d3d3d3dmZmZVVVVVVVVEREQzMzNERERmZmaIiIh3d3d3d3dmZmZVVVVVVVVERERERERVVVVVVVVVVVVVVVVERERVVVVEREREREREREREREQzMzMzMzMzMzNERERmZmZmZmZ3d3dmZmZmZmZmZmZ3d3d3d3dmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZERERERERVVVVVVVVmZmZmZmZmZmZmZmZVVVVmZmZVVVVERERVVVVVVVVVVVVERERERERERERERERERERERERERERERERERERERERVVVVmZmZmZmZmZmZmZmZVVVVVVVVERERERERERERERERVVVVVVVVERERVVVVERERERERERERERERVVVVERERVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERVVVVVVVVERERVVVVERERVVVVERERVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZ3d3dmZmZVVVVVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzNERERERERERERERERVVVVVVVUzMzMzMzMzMzMzMzMiIiIiIiIiIiJEREREREQzMzMiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIzMzMzMzMzMzMzMzNERERVVVUzMzMzMzNERERmZmZmZmZmZmZ3d3dVVVVmZmZmZmZmZmZVVVVmZmZmZmZVVVVEREREREREREREREQzMzMzMzMzMzNERERERERERERERERVVVVmZmZVVVVVVVVEREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERERERERERERERVVVVERERVVVVEREQzMzMzMzNEREQzMzN3d3d3d3dVVVVERERERERERERVVVVVVVVEREREREREREQiIiIzMzMzMzNEREQzMzMiIiIiIiIiIiIzMzMzMzNEREREREREREREREQzMzMzMzNEREQzMzMzMzNEREQzMzMzMzMzMzMzMzNEREQzMzNEREREREREREREREREREREREREREQzMzNEREREREQzMzMzMzNEREREREQzMzMzMzMzMzMzMzNERERmZmZVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERERERVVVVVVVVERERERERERERERERERERERERERERERERERERVVVVVVVUzMzNEREQzMzMzMzMzMzMzMzMiIiIzMzMzMzNVVVVmZmZmZmZEREQzMzNERERERERERERVVVVmZmZVVVVERERERERERERERERERERERERERERERERERERERERERERERERERERmZmaIiIh3d3dVVVVERERVVVVVVVVERERERERVVVVmZmZmZmZmZmZ3d3eIiIhERERERESIiIjMzMzMzMzMzMyqqqqIiIh3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERmZmZmZmZVVVVVVVVmZmZ3d3dmZmZVVVVVVVVmZmZ3d3d3d3eIiIh3d3dmZmZERERVVVVVVVVVVVVVVVVERERERERERERERERERERVVVVVVVVVVVVVVVWIiIiZmZlmZmZVVVVERERVVVVERERERERmZmaqqqqZmZlmZmZVVVVVVVWZmZmqqqqZmZmqqqqZmZl3d3dmZmZVVVV3d3eqqqqqqqqZmZmIiIiIiIiqqqqZmZmIiIh3d3dVVVVERERERERERERERERERERVVVVERERVVVVVVVVVVVVmZmZ3d3d3d3eIiIiZmZmqqqqqqqq7u7vMzMzMzMy7u7vd3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////7u7u3d3dzMzMzMzMzMzMzMzMzMzM3d3dzMzM3d3d3d3d3d3dzMzMzMzMu7u7u7u7qqqqmZmZmZmZmZmZmZmZmZmZmZmZqqqqqqqqqqqqqqqqqqqqqqqqqqqqmZmZmZmZmZmZmZmZmZmZiIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiImZmZiIiIiIiIiIiId3d3iIiIiIiIiIiIiIiIiIiImZmZmZmZmZmZmZmZiIiImZmZmZmZqqqqmZmZmZmZmZmZqqqqmZmZqqqqmZmZmZmZmZmZmZmZmZmZmZmZmZmZqqqqmZmZmZmZqqqqqqqqmZmZmZmZmZmZmZmZiIiIiIiImZmZmZmZiIiImZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZiIiImZmZmZmZmZmZmZmZiIiIiIiIiIiIiIiId3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3iIiId3d3d3d3ZmZmd3d3d3d3d3d3iIiId3d3ZmZmd3d3iIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREREREREREZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREREREVVVVREREREREREREREREREREZmZmd3d3ZmZmZmZmZmZmd3d3ZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmd3d3d3d3ZmZmZmZmd3d3d3d3d3d3d3d3ZmZmZmZmd3d3iIiIZmZmZmZmd3d3d3d3d3d3iIiIiIiIiIiId3d3ZmZmVVVVZmZmd3d3d3d3iIiIiIiIZmZmVVVVVVVVd3d3d3d3d3d3ZmZmZmZmZmZmZmZmd3d3d3d3iIiId3d3VVVVVVVVVVVVVVVVREREREREREREREREd3d3qqqqmZmZiIiIiIiId3d3ZmZmiIiIqqqqqqqqiIiId3d3d3d3d3d3ZmZmZmZmVVVVZmZmd3d3ZmZmZmZmmZmZqqqqmZmZZmZmZmZmd3d3d3d3ZmZmd3d3d3d3d3d3ZmZmVVVVREREZmZmd3d3iIiImZmZiIiId3d3d3d3d3d3d3d3iIiImZmZmZmZiIiIiIiId3d3d3d3iIiImZmZZmZmREREREREVVVVVVVVVVVVVVVVMzMzMzMzMzMzMzMzREREZmZmVVVVVVVVVVVVMzMzMzMzMzMzVVVVmZmZmZmZiIiIZmZmd3d3iIiImZmZmZmZiIiId3d3d3d3mZmZmZmZiIiId3d3ZmZmVVVVVVVVVVVVZmZmiIiId3d3ZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmVVVVVVVVVVVVVVVVZmZmd3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmVVVVREREVVVVVVVVREREREREREREREREd3d3iIiImZmZiIiIiIiIqqqqmZmZmZmZiIiIiIiId3d3d3d3d3d3d3d3d3d3iIiId3d3ZmZmd3d3qqqqmZmZiIiId3d3iIiIiIiImZmZiIiIiIiIZmZmVVVVZmZmVVVVZmZmVVVVZmZmVVVVZmZmiIiIiIiImZmZmZmZmZmZmZmZmZmZiIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiImZmZmZmZqqqqu7u7zMzMu7u7mZmZiIiIiIiIiIiId3d3ZmZmZmZmVVVVZmZmZmZmd3d3d3d3ZmZmZmZmd3d3iIiIiIiImZmZqqqqd3d3d3d3iIiImZmZd3d3ZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3VVVVVVVVVVVVd3d3iIiImZmZiIiIZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmVVVVZmZmZmZmd3d3d3d3d3d3VVVVREREZmZmd3d3d3d3iIiIiIiId3d3d3d3d3d3d3d3iIiId3d3iIiIiIiImZmZmZmZmZmZiIiIiIiId3d3d3d3d3d3iIiImZmZiIiIiIiIiIiIZmZmZmZmREREVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmVVVVVVVVREREMzMzMzMzMzMzZmZmd3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVREREREREREREREREREREREREMzMzREREREREd3d3d3d3d3d3ZmZmZmZmd3d3d3d3ZmZmd3d3ZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3ZmZmVVVVVVVVREREREREREREVVVVd3d3ZmZmZmZmVVVVZmZmZmZmVVVVVVVVZmZmVVVVREREREREREREREREREREVVVVREREMzMzREREREREVVVVREREZmZmd3d3ZmZmZmZmZmZmVVVVREREREREREREREREREREREREVVVVREREREREREREREREREREREREREREREREREREMzMzVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVREREVVVVVVVVVVVVVVVVREREVVVVREREVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVd3d3ZmZmZmZmZmZmREREREREREREREREMzMzMzMzREREVVVVREREREREREREMzMzMzMzMzMzREREREREVVVVREREMzMzIiIiMzMzMzMzIiIiMzMzMzMzREREZmZmREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzREREMzMzMzMzREREZmZmd3d3VVVVVVVVZmZmZmZmd3d3ZmZmZmZmd3d3ZmZmVVVVREREREREMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREVVVVREREVVVVREREVVVVREREREREREREREREMzMzMzMzREREVVVVmZmZiIiIVVVVREREREREREREVVVVREREREREMzMzIiIiIiIiMzMzREREMzMzIiIiIiIiMzMzMzMzREREMzMzMzMzREREMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREREREREREREREREREREREREREREREREREREREREREVVVVREREREREMzMzMzMzMzMzMzMzVVVVZmZmVVVVMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzREREVVVVZmZmVVVVVVVVVVVVd3d3ZmZmVVVVVVVVVVVVVVVVREREREREREREVVVVREREREREREREREREREREREREREREREREREREVVVVVVVVMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzREREZmZmZmZmZmZmVVVVREREREREREREVVVVVVVVVVVVREREREREVVVVREREREREMzMzREREMzMzREREMzMzREREREREREREZmZmd3d3d3d3ZmZmVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmmZmZiIiIREREVVVVu7u77u7u7u7u3d3dqqqqiIiIiIiIiIiId3d3d3d3ZmZmZmZmZmZmVVVVVVVVREREREREVVVViIiId3d3iIiIiIiIZmZmd3d3VVVVVVVVd3d3iIiIiIiId3d3ZmZmZmZmVVVVVVVVZmZmd3d3VVVVVVVVVVVVVVVVREREREREVVVVVVVVVVVVVVVVVVVViIiIzMzMqqqqd3d3VVVVVVVVREREREREZmZmmZmZu7u7iIiIVVVVVVVVmZmZu7u7mZmZqqqqmZmZiIiId3d3ZmZmd3d3mZmZmZmZiIiIiIiImZmZmZmZiIiImZmZmZmZZmZmVVVVREREREREREREREREVVVVREREVVVVVVVVREREVVVVZmZmd3d3d3d3d3d3iIiIqqqqqqqqqqqqzMzMu7u7zMzM3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////+7u7t3d3d3d3e7u7t3d3e7u7u7u7u7u7t3d3e7u7t3d3e7u7u7u7t3d3d3d3czMzMzMzLu7u6qqqqqqqru7u6qqqqqqqru7u7u7u8zMzMzMzMzMzMzMzMzMzLu7u8zMzMzMzMzMzMzMzLu7u7u7u6qqqqqqqpmZmZmZmZmZmZmZmZmZmZmZmYiIiJmZmZmZmaqqqqqqqru7u7u7u7u7u7u7u7u7u7u7u6qqqqqqqru7u6qqqru7u6qqqqqqqqqqqqqqqqqqqqqqqpmZmZmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d2ZmZmZmZlVVVVVVVWZmZlVVVWZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZnd3d2ZmZmZmZnd3d3d3d3d3d4iIiHd3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d2ZmZmZmZnd3d2ZmZmZmZnd3d3d3d4iIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiHd3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVURERERERERERERERDMzM0RERFVVVWZmZnd3d2ZmZlVVVWZmZmZmZmZmZmZmZlVVVVVVVXd3d2ZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZoiIiHd3d2ZmZmZmZnd3d4iIiIiIiIiIiIiIiIiIiHd3d2ZmZmZmZmZmZoiIiHd3d3d3d3d3d3d3d2ZmZnd3d4iIiJmZmXd3d2ZmZmZmZmZmZmZmZmZmZnd3d6qqqoiIiFVVVVVVVURERERERFVVVURERFVVVWZmZpmZmczMzLu7u6qqqpmZmXd3d4iIiKqqqru7u7u7u6qqqpmZmZmZmYiIiHd3d4iIiHd3d2ZmZmZmZoiIiJmZmaqqqqqqqqqqqoiIiIiIiIiIiHd3d3d3d4iIiIiIiHd3d2ZmZnd3d2ZmZnd3d3d3d4iIiJmZmZmZmZmZmZmZmZmZmZmZmZmZmbu7u6qqqpmZmZmZmYiIiHd3d6qqqru7u2ZmZkRERDMzM2ZmZlVVVVVVVWZmZkRERDMzMzMzMzMzMzMzM1VVVVVVVWZmZmZmZkRERDMzMzMzM2ZmZqqqqqqqqoiIiHd3d3d3d2ZmZpmZmZmZmZmZmYiIiHd3d3d3d4iIiIiIiHd3d2ZmZmZmZkRERDMzM0RERIiIiJmZmXd3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZlVVVVVVVWZmZlVVVVVVVWZmZnd3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZlVVVWZmZmZmZkRERERERERERFVVVVVVVXd3d4iIiIiIiJmZmYiIiIiIiIiIiJmZmYiIiIiIiHd3d3d3d2ZmZmZmZnd3d3d3d2ZmZnd3d5mZmaqqqqqqqpmZmZmZmZmZmaqqqpmZmXd3d2ZmZlVVVWZmZnd3d2ZmZmZmZmZmZnd3d3d3d2ZmZoiIiKqqqpmZmYiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d4iIiHd3d3d3d3d3d4iIiJmZmZmZmZmZmaqqqru7u7u7u6qqqoiIiHd3d3d3d3d3d1VVVVVVVWZmZmZmZmZmZmZmZnd3d4iIiGZmZnd3d3d3d3d3d2ZmZmZmZoiIiIiIiJmZmYiIiHd3d1VVVVVVVWZmZlVVVVVVVVVVVVVVVWZmZmZmZnd3d4iIiHd3d2ZmZlVVVWZmZoiIiKqqqpmZmYiIiHd3d3d3d2ZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZlVVVWZmZnd3d3d3d5mZmYiIiHd3d4iIiIiIiIiIiIiIiHd3d4iIiJmZmZmZmZmZmZmZmYiIiIiIiIiIiIiIiHd3d3d3d5mZmZmZmYiIiIiIiHd3d1VVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVURERERERFVVVURERDMzMzMzMzMzM1VVVXd3d3d3d4iIiHd3d2ZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVURERERERDMzMzMzMzMzM2ZmZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZnd3d2ZmZnd3d3d3d3d3d2ZmZmZmZnd3d3d3d2ZmZlVVVURERFVVVVVVVURERGZmZnd3d2ZmZmZmZmZmZlVVVVVVVWZmZlVVVVVVVURERERERERERERERERERFVVVURERERERERERERERERERERERERERGZmZnd3d3d3d2ZmZmZmZlVVVURERERERDMzMzMzMzMzMzMzM0RERERERDMzMzMzMzMzM0RERDMzMzMzMzMzM0RERERERFVVVWZmZkRERGZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVURERFVVVWZmZmZmZmZmZmZmZlVVVURERERERERERDMzM0RERERERFVVVURERERERERERDMzMzMzMzMzMzMzM0RERERERERERDMzMyIiIiIiIjMzMzMzMyIiIkRERERERFVVVURERDMzMyIiIjMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzM0RERDMzMzMzM0RERERERFVVVWZmZlVVVVVVVVVVVWZmZnd3d4iIiHd3d3d3d1VVVURERERERDMzM0RERDMzM0RERERERERERERERDMzMzMzM0RERERERERERFVVVURERERERERERDMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVURERFVVVVVVVURERERERFVVVURERERERDMzM1VVVXd3d5mZmXd3d0RERERERERERERERDMzM0RERDMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIiIiIjMzM0RERERERDMzM0RERDMzM0RERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzM0RERDMzM0RERERERERERERERERERERERERERDMzMzMzM1VVVVVVVVVVVURERGZmZlVVVURERDMzMzMzM1VVVWZmZlVVVURERDMzMzMzMzMzMzMzM0RERDMzM0RERERERDMzM1VVVVVVVWZmZlVVVVVVVVVVVWZmZnd3d3d3d2ZmZmZmZlVVVURERERERFVVVURERERERERERERERERERERERERERERERERERERERFVVVWZmZlVVVTMzM0RERDMzM0RERDMzM0RERERERDMzM0RERGZmZmZmZmZmZkRERERERERERFVVVVVVVVVVVURERERERERERERERERERERERERERDMzM0RERDMzM0RERDMzM0RERERERHd3d3d3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d2ZmZmZmZnd3d3d3dzMzM2ZmZt3d3e7u7u7u7u7u7ru7u5mZmYiIiIiIiIiIiIiIiHd3d2ZmZmZmZlVVVVVVVURERFVVVWZmZpmZmXd3d2ZmZnd3d2ZmZlVVVVVVVWZmZoiIiIiIiGZmZlVVVVVVVWZmZlVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVaqqqszMzIiIiFVVVURERFVVVVVVVURERFVVVZmZmZmZmVVVVURERHd3d7u7u6qqqru7u6qqqqqqqoiIiHd3d3d3d4iIiIiIiIiIiJmZmZmZmYiIiHd3d3d3d3d3d3d3d3d3d1VVVURERERERFVVVVVVVURERFVVVURERERERERERFVVVVVVVXd3d4iIiHd3d5mZmZmZmZmZmaqqqru7u8zMzMzMzN3d3d3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////u7u7u7u7d3d3d3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMy7u7u7u7u7u7vMzMy7u7u7u7uqqqq7u7u7u7u7u7u7u7vMzMzMzMzd3d3d3d3MzMzd3d3MzMzd3d3MzMzMzMzMzMy7u7vMzMzMzMzMzMy7u7u7u7uqqqq7u7u7u7u7u7u7u7vMzMzMzMzMzMzd3d3d3d3MzMzMzMzMzMzMzMzMzMzMzMzd3d3MzMzMzMzMzMzMzMy7u7vMzMy7u7u7u7uqqqqqqqqZmZmZmZmqqqqZmZmqqqqZmZmqqqqZmZmZmZmIiIiIiIiIiIh3d3dVVVVVVVVERERERERERERERERERERERERERERERERERERERERVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3eIiIiIiIiIiIiIiIiZmZmZmZmIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIh3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVEREREREQzMzNEREQzMzMzMzMzMzMzMzNmZmZ3d3dmZmZERERmZmZmZmZmZmZmZmZVVVVmZmZ3d3dmZmZVVVV3d3dmZmZVVVVmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZ3d3eIiIh3d3eIiIiIiIiIiIiIiIiZmZmZmZmIiIh3d3dmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIiqqqqZmZlmZmZVVVVmZmZmZmZVVVVmZmaIiIiZmZl3d3dVVVVVVVVVVVVVVVVERERVVVVVVVV3d3eqqqrd3d3MzMzMzMyqqqqZmZmZmZm7u7u7u7uqqqqqqqqqqqqqqqqqqqqIiIiZmZmZmZl3d3d3d3eZmZmqqqqqqqqqqqqqqqqqqqqqqqqZmZmIiIiIiIiIiIiIiIh3d3eIiIh3d3eIiIiZmZmIiIiIiIiIiIiZmZmqqqqqqqqqqqqqqqqZmZm7u7u7u7uqqqqIiIiIiIh3d3eIiIi7u7uIiIhERERERERERERVVVVVVVVmZmZEREQzMzNERERERERERERVVVVVVVVVVVVEREREREQzMzNERERmZmaZmZmqqqqZmZmIiIhmZmaIiIiZmZmZmZmIiIh3d3d3d3d3d3eIiIiIiIhmZmZmZmZVVVVERERERERERER3d3eZmZl3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3dmZmZ3d3dmZmZmZmZVVVVVVVVERERVVVV3d3eIiIh3d3dmZmZ3d3d3d3d3d3d3d3dmZmZmZmZmZmZERERVVVVVVVUzMzNERERVVVVVVVVVVVVmZmaIiIiZmZmIiIiIiIiIiIiIiIiIiIiZmZmIiIh3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmaZmZmqqqq7u7u7u7u7u7u7u7uZmZmIiIh3d3dmZmZmZmZ3d3d3d3dmZmZmZmZVVVVmZmZ3d3d3d3eIiIiqqqqZmZmZmZmIiIh3d3eIiIiIiIiZmZl3d3d3d3eIiIiIiIh3d3d3d3d3d3d3d3eIiIiZmZl3d3eIiIiZmZmqqqqqqqqIiIiIiIh3d3dmZmZVVVVmZmZ3d3dmZmZmZmZmZmZ3d3eIiIh3d3d3d3dmZmZVVVVmZmZVVVV3d3eZmZmZmZmZmZl3d3dmZmZVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZ3d3eIiIiIiIh3d3dVVVVmZmaZmZmqqqqZmZmZmZl3d3d3d3d3d3d3d3d3d3d3d3dmZmaIiIh3d3dmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZ3d3eZmZmIiIiIiIiIiIiIiIiIiIh3d3eIiIiZmZmZmZmZmZmIiIiIiIiZmZl3d3eIiIiZmZl3d3dmZmaZmZmZmZmZmZl3d3dmZmZmZmZVVVVVVVVmZmZVVVVVVVVERERVVVVERERERERVVVVEREREREQzMzMiIiIzMzNVVVVmZmaIiIiIiIh3d3d3d3dmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVVERERERERERERERERVVVVEREQzMzMzMzMzMzNmZmZ3d3d3d3d3d3d3d3dmZmZmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZ3d3dmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVERERVVVVVVVVERERERERERERVVVUzMzMzMzNERERERERERERERERVVVV3d3dmZmZmZmZmZmZVVVVVVVVEREREREQzMzNEREQzMzNEREREREQzMzMzMzMzMzNEREQzMzMzMzMzMzNERERERERVVVVmZmZVVVVmZmZ3d3dmZmZVVVVVVVVVVVVVVVVERERVVVVmZmZVVVVVVVVVVVVERERERERERERERERERERERERERERERERVVVVVVVVVVVV3d3dmZmZ3d3dVVVVEREREREREREQzMzMzMzMzMzNERERVVVUzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMiIiIiIiIzMzMzMzMiIiIzMzNEREREREREREQzMzMiIiIiIiIiIiIiIiIzMzMzMzMzMzMiIiIiIiIREREiIiIiIiIzMzNERERVVVVEREREREREREQzMzNVVVVERERVVVVVVVVVVVVmZmZmZmZ3d3eIiIh3d3dmZmZVVVVEREREREQzMzMzMzNEREREREREREREREQzMzMzMzMzMzNEREQzMzNERERERERVVVVVVVVEREREREQzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERVVVVVVVVVVVVVVVVERERERERVVVVEREQzMzMzMzNERERVVVWIiIiZmZlmZmZEREREREREREREREQzMzNEREQzMzMzMzMiIiIiIiIzMzMzMzMiIiIiIiIzMzMzMzNEREREREQzMzNEREQzMzNEREREREREREQzMzMzMzMzMzNEREQzMzNEREREREQzMzNEREREREQzMzNEREREREREREREREREREREREREREQzMzNERERERERmZmZVVVVERERERERmZmZVVVVEREQzMzMiIiJERERVVVVEREREREREREQzMzNEREREREREREREREQzMzNERERERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZVVVVERERERERVVVVVVVVEREREREREREREREREREREREREREREREQzMzNERERVVVVVVVVEREQzMzMzMzNEREQzMzNEREREREQzMzNERERVVVVmZmZVVVVVVVVVVVVERERERERVVVV3d3dmZmZERERERERERERERERVVVVEREQzMzNEREREREQzMzNEREQzMzNERERVVVV3d3dmZmZVVVVVVVVVVVVERERVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVV3d3dmZmZERER3d3fd3d3////u7u7u7u7MzMyZmZmZmZmIiIiIiIiIiIh3d3d3d3dmZmZmZmZVVVVERERVVVVmZmZ3d3dmZmZmZmZmZmZVVVVVVVVVVVVVVVV3d3d3d3dmZmZVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVmZmZVVVVmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVVVVWIiIi7u7uIiIhVVVVVVVVVVVVERERERERVVVWZmZmqqqpmZmYzMzN3d3eqqqq7u7u7u7uqqqqqqqqZmZmIiIh3d3dmZmZ3d3eIiIiIiIiIiIiZmZmIiIhmZmZVVVWIiIiZmZlmZmZEREQzMzNVVVVERERERERERERVVVVVVVVERERERERVVVVmZmaIiIiIiIiIiIiZmZmIiIiZmZmqqqq7u7vMzMzMzMzd3d3u7u7u7u7////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////7u7u////////////////////////7u7u3d3d3d3d3d3dzMzM3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM3d3dzMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7u7u7zMzMzMzM3d3d3d3d3d3d3d3d3d3d7u7u3d3d3d3d3d3dzMzMzMzMzMzM3d3dzMzM3d3dzMzMzMzMu7u7zMzMzMzMzMzMzMzMzMzMzMzMzMzM3d3dzMzM3d3dzMzMzMzMzMzM3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzM3d3dzMzMzMzMu7u7zMzMu7u7u7u7zMzMu7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqmZmZiIiId3d3VVVVVVVVREREREREMzMzREREMzMzREREMzMzMzMzREREREREREREMzMzREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3iIiIiIiIiIiIiIiIiIiImZmZiIiIiIiIiIiIiIiIiIiImZmZiIiImZmZiIiIiIiIiIiId3d3iIiIiIiIiIiImZmZiIiIiIiIiIiIiIiIiIiIiIiId3d3ZmZmVVVVZmZmVVVVVVVVVVVVVVVVREREMzMzMzMzMzMzMzMzVVVVZmZmZmZmREREREREZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmd3d3VVVVVVVVZmZmZmZmZmZmd3d3d3d3ZmZmd3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIZmZmZmZmZmZmd3d3d3d3iIiIiIiId3d3iIiIiIiImZmZqqqqiIiId3d3ZmZmZmZmZmZmVVVVZmZmd3d3d3d3d3d3ZmZmZmZmVVVVVVVVMzMzREREd3d3iIiIqqqqzMzM3d3dzMzMu7u7u7u7zMzMzMzMu7u7qqqqmZmZqqqqu7u7u7u7iIiIiIiImZmZiIiImZmZzMzM3d3du7u7qqqqu7u7qqqqmZmZmZmZiIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3iIiImZmZmZmZmZmZmZmZiIiImZmZmZmZmZmZqqqqqqqqqqqqmZmZmZmZiIiId3d3d3d3mZmZiIiIREREMzMzVVVVREREVVVVVVVVREREMzMzREREZmZmVVVVVVVVREREMzMzREREMzMzVVVVVVVVREREd3d3mZmZu7u7qqqqiIiId3d3iIiImZmZqqqqiIiIZmZmZmZmiIiIiIiIZmZmVVVVVVVVVVVVREREREREd3d3mZmZiIiIiIiIiIiId3d3d3d3d3d3iIiIiIiId3d3d3d3d3d3ZmZmVVVVZmZmVVVVVVVVREREZmZmmZmZqqqqiIiIiIiIiIiId3d3ZmZmVVVVVVVVVVVVVVVVREREREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3iIiIiIiId3d3iIiId3d3iIiId3d3iIiIiIiId3d3ZmZmZmZmZmZmZmZmd3d3ZmZmiIiIqqqqqqqqu7u7qqqqmZmZd3d3d3d3ZmZmZmZmZmZmVVVVZmZmVVVVVVVVZmZmZmZmd3d3d3d3iIiImZmZmZmZiIiId3d3iIiImZmZiIiId3d3iIiIiIiIiIiImZmZiIiIiIiId3d3iIiIiIiIiIiId3d3d3d3iIiIqqqqmZmZiIiId3d3d3d3VVVVZmZmd3d3ZmZmVVVVZmZmZmZmd3d3iIiId3d3ZmZmVVVVZmZmZmZmd3d3mZmZmZmZiIiIZmZmVVVVVVVVZmZmZmZmZmZmd3d3ZmZmVVVVZmZmZmZmd3d3d3d3d3d3ZmZmZmZmqqqqu7u7qqqqiIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3iIiId3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmd3d3iIiIiIiImZmZiIiIiIiImZmZmZmZiIiIiIiIiIiIiIiImZmZmZmZmZmZiIiIiIiIiIiIiIiIZmZmVVVViIiIiIiImZmZiIiIZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVREREREREREREREREREREREREMzMzMzMzMzMzVVVVZmZmd3d3iIiId3d3d3d3ZmZmVVVVZmZmVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREMzMzMzMzMzMzVVVVd3d3d3d3iIiIZmZmd3d3d3d3ZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVZmZmd3d3d3d3ZmZmd3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREMzMzMzMzREREREREMzMzMzMzREREREREREREREREREREVVVVZmZmZmZmZmZmZmZmREREREREMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzREREREREREREMzMzREREMzMzREREREREZmZmVVVVZmZmZmZmZmZmVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVREREVVVVREREVVVVREREREREREREREREREREREREVVVVZmZmZmZmZmZmZmZmZmZmVVVVREREREREMzMzMzMzMzMzREREREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzMzMzMzMzREREREREMzMzMzMzIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzREREVVVVREREREREREREMzMzMzMzREREREREREREREREVVVVZmZmZmZmZmZmZmZmZmZmVVVVREREMzMzREREMzMzREREREREVVVVREREREREREREMzMzMzMzREREREREMzMzREREREREREREREREREREREREREREREREREREREREMzMzMzMzREREMzMzREREMzMzMzMzMzMzREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREMzMzREREVVVVd3d3iIiIZmZmREREVVVVREREREREMzMzMzMzMzMzIiIiIiIiMzMzREREMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREMzMzREREMzMzREREMzMzREREMzMzMzMzMzMzREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREVVVVZmZmVVVVREREREREVVVVVVVVVVVVREREMzMzREREVVVVREREMzMzMzMzREREREREREREMzMzREREREREMzMzREREREREVVVVVVVVREREREREVVVVZmZmVVVVREREVVVVREREVVVVREREREREVVVVREREVVVVREREREREREREREREREREMzMzREREREREREREVVVVREREREREMzMzREREREREMzMzREREMzMzREREREREVVVVVVVVZmZmZmZmREREREREVVVVd3d3ZmZmVVVVREREREREVVVVREREREREREREREREREREMzMzREREMzMzVVVVZmZmZmZmVVVVVVVVZmZmVVVVVVVVVVVVREREVVVVZmZmZmZmZmZmd3d3ZmZmd3d3d3d3REREd3d33d3d7u7u7u7u7u7uzMzMqqqqiIiIiIiImZmZiIiIiIiIiIiIZmZmVVVVVVVVVVVVVVVVZmZmVVVVZmZmd3d3d3d3VVVVVVVVREREVVVVVVVVVVVVZmZmZmZmREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVREREREREREREVVVVVVVVZmZmiIiImZmZd3d3VVVVVVVVVVVVREREVVVVmZmZu7u7ZmZmMzMzZmZmu7u7zMzMu7u7qqqqu7u7u7u7mZmZiIiId3d3iIiIiIiImZmZu7u7zMzMu7u7mZmZZmZmiIiIqqqqiIiIVVVVREREREREREREREREREREREREVVVVREREVVVVREREVVVVZmZmiIiIiIiIiIiIiIiId3d3iIiImZmZu7u7u7u7zMzMzMzM7u7u7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////+7u7v///////////+7u7u7u7t3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzN3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzN3d3d3d3d3d3czMzMzMzN3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3czMzMzMzMzMzN3d3czMzN3d3czMzN3d3czMzMzMzN3d3czMzN3d3czMzMzMzMzMzLu7u8zMzMzMzLu7u7u7u7u7u5mZmZmZmYiIiHd3d2ZmZlVVVVVVVVVVVURERFVVVURERERERERERERERERERDMzM0RERDMzM0RERDMzM0RERDMzMzMzMzMzM0RERERERERERERERERERERERERERERERERERFVVVURERFVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d4iIiIiIiJmZmYiIiIiIiIiIiJmZmYiIiIiIiJmZmYiIiIiIiJmZmZmZmZmZmZmZmYiIiIiIiIiIiIiIiHd3d2ZmZmZmZmZmZkRERFVVVVVVVURERERERERERDMzM1VVVVVVVURERFVVVVVVVWZmZmZmZmZmZnd3d3d3d2ZmZmZmZmZmZlVVVVVVVWZmZnd3d2ZmZoiIiJmZmYiIiIiIiIiIiIiIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d2ZmZnd3d3d3d3d3d4iIiJmZmYiIiIiIiJmZmYiIiIiIiIiIiHd3d3d3d3d3d2ZmZlVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZkRERERERERERERERGZmZpmZmaqqqru7u8zMzKqqqru7u8zMzN3d3d3d3czMzLu7u6qqqru7u7u7u7u7u6qqqpmZmYiIiHd3d7u7u93d3d3d3czMzLu7u7u7u6qqqpmZmaqqqqqqqoiIiHd3d3d3d4iIiGZmZnd3d3d3d4iIiKqqqqqqqpmZmYiIiIiIiJmZmZmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiIiIiHd3d3d3d2ZmZjMzM0RERHd3d3d3d3d3d2ZmZkRERERERERERGZmZmZmZkRERERERDMzMyIiIjMzM1VVVVVVVURERFVVVZmZmbu7u6qqqoiIiIiIiIiIiJmZmaqqqpmZmWZmZnd3d3d3d3d3d3d3d2ZmZmZmZkRERERERFVVVXd3d5mZmZmZmYiIiHd3d3d3d4iIiIiIiJmZmYiIiHd3d1VVVVVVVWZmZmZmZlVVVVVVVWZmZlVVVVVVVYiIiLu7u6qqqoiIiHd3d3d3d3d3d1VVVURERFVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVXd3d2ZmZnd3d5mZmYiIiHd3d3d3d2ZmZmZmZnd3d3d3d3d3d2ZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d5mZmaqqqpmZmXd3d2ZmZnd3d2ZmZlVVVWZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZoiIiGZmZmZmZnd3d3d3d4iIiIiIiIiIiHd3d4iIiIiIiIiIiJmZmZmZmaqqqoiIiJmZmZmZmZmZmYiIiHd3d2ZmZmZmZoiIiJmZmXd3d3d3d2ZmZlVVVWZmZlVVVWZmZnd3d2ZmZmZmZnd3d4iIiHd3d3d3d2ZmZnd3d2ZmZoiIiJmZmXd3d3d3d2ZmZmZmZlVVVWZmZlVVVWZmZmZmZlVVVVVVVXd3d3d3d2ZmZmZmZnd3d2ZmZlVVVZmZmbu7u6qqqpmZmYiIiHd3d3d3d3d3d3d3d2ZmZnd3d3d3d3d3d4iIiIiIiHd3d3d3d3d3d3d3d4iIiJmZmYiIiIiIiIiIiJmZmYiIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d0RERGZmZpmZmZmZmYiIiIiIiHd3d2ZmZlVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVURERERERDMzMzMzMzMzM1VVVVVVVWZmZnd3d4iIiGZmZlVVVVVVVWZmZmZmZlVVVWZmZmZmZlVVVVVVVURERFVVVVVVVVVVVURERERERFVVVVVVVVVVVXd3d4iIiGZmZnd3d3d3d2ZmZmZmZmZmZmZmZnd3d1VVVVVVVWZmZlVVVVVVVWZmZmZmZlVVVWZmZmZmZlVVVVVVVVVVVWZmZnd3d2ZmZmZmZlVVVURERERERFVVVVVVVVVVVURERDMzMzMzMzMzMzMzM0RERERERDMzMzMzM0RERFVVVWZmZlVVVURERFVVVWZmZmZmZmZmZkRERERERDMzM0RERERERDMzMzMzM0RERDMzM0RERERERDMzMzMzMzMzM0RERERERERERERERFVVVWZmZnd3d2ZmZlVVVVVVVVVVVURERERERFVVVVVVVURERERERERERERERERERERERERERFVVVURERERERDMzM0RERERERFVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERERERERERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIjMzM0RERERERERERERERERERERERDMzMzMzM0RERDMzM0RERERERFVVVVVVVVVVVWZmZlVVVVVVVURERERERERERERERERERERERFVVVTMzMzMzM0RERDMzMzMzMzMzM0RERERERERERERERERERERERERERERERERERERERERERDMzM0RERDMzMzMzMzMzM0RERDMzMzMzMzMzMzMzM0RERFVVVVVVVURERFVVVWZmZlVVVWZmZlVVVURERERERERERERERHd3d4iIiGZmZlVVVURERERERERERERERDMzMzMzMzMzMyIiIjMzM0RERERERDMzMzMzMzMzM0RERDMzM0RERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERDMzM0RERERERERERERERERERDMzM0RERERERERERERERERERERERGZmZmZmZlVVVURERERERERERERERFVVVVVVVTMzM0RERFVVVTMzMzMzMzMzMzMzM0RERERERERERDMzMzMzM0RERERERDMzM0RERERERERERERERFVVVVVVVVVVVURERFVVVVVVVVVVVURERERERERERERERERERERERERERERERERERERERDMzMzMzM0RERGZmZkRERDMzMzMzM0RERFVVVVVVVURERERERERERFVVVVVVVVVVVVVVVYiIiIiIiERERDMzM1VVVXd3d2ZmZkRERERERERERERERFVVVVVVVURERERERERERERERERERFVVVWZmZnd3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVXd3d3d3d3d3d2ZmZnd3d3d3d0RERHd3d93d3d3d3e7u7t3d3bu7u5mZmYiIiIiIiJmZmYiIiJmZmXd3d3d3d2ZmZlVVVWZmZnd3d2ZmZlVVVVVVVXd3d4iIiGZmZkRERFVVVVVVVVVVVVVVVVVVVVVVVURERERERERERGZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVVVVVURERFVVVURERFVVVVVVVVVVVVVVVZmZmczMzHd3d1VVVVVVVURERERERFVVVYiIiLu7u3d3d0RERGZmZqqqqru7u7u7u6qqqru7u7u7u4iIiIiIiHd3d2ZmZnd3d6qqqru7u7u7u7u7u5mZmYiIiJmZmZmZmYiIiIiIiHd3d1VVVVVVVURERERERFVVVURERERERERERERERERERFVVVXd3d5mZmYiIiHd3d4iIiHd3d5mZmZmZmaqqqru7u7u7u8zMzN3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////u7u7d3d3MzMy7u7u7u7u7u7vMzMzMzMy7u7u7u7vMzMzMzMzd3d3MzMzd3d3d3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3MzMzMzMy7u7vMzMy7u7u7u7u7u7u7u7u7u7uqqqq7u7u7u7u7u7u7u7u7u7u7u7u7u7vMzMzMzMzMzMzd3d3d3d3u7u7d3d3d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzd3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3MzMzMzMzMzMy7u7vMzMy7u7u7u7u7u7u7u7uqqqqqqqqZmZmZmZmIiIiIiIh3d3d3d3dmZmZ3d3dmZmZmZmZVVVVmZmZVVVVVVVVEREREREREREREREREREREREREREQzMzNEREREREREREQzMzNEREQzMzMzMzNERERERERERERERERERERERERERERERERVVVVERERVVVVVVVVVVVVVVVVVVVV3d3dmZmZ3d3d3d3eIiIh3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZVVVVVVVVVVVVmZmZmZmZ3d3eZmZmZmZmqqqqZmZmIiIiIiIiIiIh3d3d3d3d3d3dmZmZ3d3d3d3eIiIiIiIiIiIiIiIh3d3d3d3eIiIh3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3dmZmZ3d3dmZmZVVVVmZmZ3d3dmZmZVVVVVVVVVVVVERERVVVVERERERERmZmaZmZmqqqqqqqq7u7uqqqq7u7vd3d3d3d3d3d3MzMzMzMzMzMzMzMy7u7uZmZmqqqqqqqp3d3d3d3fMzMzd3d3MzMzMzMy7u7u7u7uqqqqqqqqqqqqZmZmIiIh3d3dmZmaIiIh3d3d3d3eIiIiIiIiZmZmqqqqZmZmZmZmZmZmZmZmZmZmIiIiIiIiZmZmIiIh3d3d3d3d3d3eIiIiIiIhVVVVERERERERERER3d3eIiIiIiIh3d3dEREREREREREREREREREREREREREREREQzMzMzMzNVVVVVVVVVVVVVVVV3d3eqqqqqqqqZmZmZmZmZmZmZmZmZmZmqqqqIiIh3d3d3d3d3d3dmZmZmZmZVVVVERERVVVVVVVVmZmZ3d3eZmZmZmZl3d3d3d3d3d3eZmZmIiIiIiIh3d3dmZmZmZmZmZmZmZmZVVVVVVVVmZmZVVVUzMzNVVVWZmZm7u7uIiIiIiIiIiIhmZmZmZmZEREQzMzNERERVVVVmZmZVVVVVVVVVVVVVVVVmZmZ3d3d3d3dmZmaZmZmZmZl3d3d3d3dmZmZ3d3d3d3dmZmZ3d3dmZmZ3d3d3d3dmZmZ3d3d3d3dmZmZmZmZmZmZ3d3eZmZmZmZl3d3d3d3d3d3d3d3dmZmZVVVVmZmZmZmZmZmZVVVVmZmZmZmZ3d3d3d3d3d3dVVVVVVVV3d3eIiIiZmZmIiIiIiIiZmZmqqqqZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmIiIhmZmZ3d3eIiIh3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZ3d3d3d3eIiIh3d3dmZmZmZmZ3d3eIiIiZmZmZmZlmZmZmZmZmZmZmZmZmZmZVVVVmZmZ3d3dmZmZmZmZ3d3dmZmZmZmZVVVV3d3dmZmZVVVWZmZnMzMyqqqqIiIiIiIh3d3d3d3d3d3eIiIh3d3eIiIiIiIiIiIiZmZmZmZmIiIh3d3d3d3dmZmZ3d3eqqqqZmZmIiIiIiIiIiIiIiIiIiIh3d3eIiIiIiIh3d3eIiIiZmZmIiIiIiIiIiIiIiIiIiIh3d3d3d3dVVVVVVVV3d3d3d3eIiIiIiIhVVVVVVVVVVVVVVVVERERVVVVVVVVmZmZERERVVVVVVVVEREREREREREQzMzMzMzMzMzNERERVVVVmZmaIiIiIiIh3d3dVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVERERVVVVERERVVVVERERVVVVVVVVVVVVmZmZmZmaIiIiIiIhmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVERERVVVVERERVVVVmZmZmZmZmZmZVVVVERERVVVVEREREREREREREREREREREREREREQzMzNERERVVVVEREQzMzNERERVVVVVVVVVVVVERERVVVVVVVVmZmZmZmZEREREREREREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMiIiJERERERERERERERERERERERERVVVVmZmZmZmZmZmZmZmZmZmZERERERERVVVVVVVVERERERERERERERERERERERERERERERERERERERERERERERERVVVVERERVVVVERERVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVEREREREQzMzNEREQzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIzMzMzMzMzMzMiIiIiIiIzMzNEREQzMzMzMzMzMzMzMzNERERERERERERVVVVEREREREREREQzMzMzMzNEREREREREREQzMzNERERVVVVVVVVmZmZVVVVVVVVEREREREREREREREREREREREREREREREQzMzMzMzNEREREREQzMzNEREREREREREQzMzNEREQzMzNERERVVVVVVVVVVVVEREREREREREQzMzNEREQzMzMzMzNEREQzMzMzMzMzMzNERERVVVVERERVVVVERERmZmZVVVVVVVVVVVVERERERERERERVVVV3d3d3d3dmZmZVVVVVVVVEREQzMzNEREREREQzMzMiIiIiIiJERERVVVUzMzNEREQzMzMzMzMzMzNEREREREQzMzNEREQzMzNEREQzMzMzMzMzMzNEREQzMzMzMzMzMzNERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERVVVVVVVVVVVVEREREREQzMzMzMzMzMzNERERERERVVVVmZmZEREQzMzMzMzNEREQzMzNEREREREQzMzNEREREREQzMzNERERERERERERERERERERERERVVVVVVVVERERERERVVVVVVVVEREREREREREREREREREQzMzNERERERERERERERERERERERERERER3d3dmZmYzMzMzMzNERERVVVVVVVVERERERERVVVVVVVVVVVVVVVVmZmaIiIiZmZlVVVUzMzNERERVVVV3d3dVVVVERERERERERERERERERERERERERERVVVVERERERERERERmZmZ3d3dVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZ3d3dmZmZmZmZ3d3d3d3dERERmZmaqqqrd3d3d3d3u7u7d3d2ZmZmIiIiIiIiIiIiIiIiIiIh3d3dmZmZmZmZVVVVmZmZmZmZVVVVVVVVVVVV3d3eIiIhmZmZERERVVVVVVVVVVVVVVVVVVVVERERERERERERVVVVVVVVVVVVmZmZVVVVmZmZmZmZVVVVVVVVVVVVVVVVERERERERVVVVVVVVERERVVVWZmZnMzMyIiIhVVVVVVVVVVVVERERVVVWIiIjMzMyZmZlERERmZmaqqqq7u7vMzMyqqqqqqqqZmZmIiIiIiIiIiIhmZmZmZmaIiIiqqqqZmZmqqqqZmZmIiIiqqqqZmZlVVVV3d3eqqqqIiIhmZmZmZmZVVVVVVVVERERERERERERERERERERERERVVVV3d3eZmZmIiIiIiIiIiIiIiIiIiIiZmZm7u7u7u7uZmZmZmZnMzMzu7u7u7u7////////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////7u7u////3d3du7u7u7u7u7u7u7u7zMzMzMzMzMzM3d3dzMzM3d3dzMzMzMzM3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMu7u7u7u7qqqqu7u7qqqqqqqqqqqqqqqqu7u7u7u7u7u7u7u7zMzMzMzMzMzMzMzM3d3dzMzM3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM3d3dzMzM3d3dzMzMzMzMzMzMzMzMzMzMu7u7u7u7zMzMu7u7qqqqqqqqu7u7qqqqu7u7qqqqqqqqmZmZmZmZmZmZmZmZmZmZiIiIiIiIiIiIiIiIiIiIZmZmZmZmZmZmVVVVVVVVVVVVREREVVVVREREREREREREMzMzREREMzMzMzMzMzMzREREMzMzREREMzMzREREMzMzREREREREREREREREREREREREMzMzREREVVVVREREREREVVVVVVVVVVVVZmZmd3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3iIiId3d3d3d3ZmZmVVVVZmZmVVVVVVVVREREREREVVVVVVVVREREVVVVREREREREVVVVREREREREVVVVd3d3VVVVZmZmiIiIiIiImZmZqqqqmZmZiIiIqqqqmZmZZmZmd3d3d3d3d3d3d3d3iIiImZmZmZmZmZmZiIiId3d3d3d3iIiId3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmVVVVd3d3ZmZmZmZmVVVVVVVVREREMzMzREREMzMzVVVVZmZmiIiIqqqqqqqqmZmZiIiIqqqqzMzM7u7u3d3dzMzM3d3d3d3dzMzMu7u7mZmZmZmZmZmZiIiImZmZu7u73d3d3d3dzMzMzMzMqqqqqqqqqqqqqqqqmZmZd3d3d3d3iIiIiIiId3d3ZmZmd3d3iIiImZmZmZmZqqqqmZmZiIiIiIiIiIiIiIiImZmZmZmZiIiId3d3d3d3iIiIiIiIZmZmREREMzMzREREMzMzVVVVd3d3iIiIZmZmVVVVREREVVVVREREREREMzMzMzMzMzMzMzMzMzMzREREVVVVVVVVREREVVVViIiIqqqqmZmZmZmZqqqqmZmZqqqqqqqqmZmZd3d3ZmZmd3d3VVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmiIiIiIiIiIiIiIiId3d3iIiIiIiId3d3d3d3VVVVZmZmZmZmVVVVVVVVVVVVVVVVZmZmREREREREd3d3u7u7qqqqd3d3d3d3ZmZmZmZmREREREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmd3d3d3d3ZmZmd3d3mZmZmZmZiIiId3d3d3d3d3d3ZmZmd3d3d3d3ZmZmd3d3ZmZmd3d3d3d3ZmZmZmZmZmZmZmZmd3d3d3d3iIiId3d3iIiId3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmd3d3d3d3iIiId3d3ZmZmREREd3d3mZmZqqqqmZmZiIiImZmZqqqqqqqqmZmZmZmZmZmZmZmZmZmZqqqqmZmZmZmZiIiId3d3d3d3iIiId3d3ZmZmd3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3ZmZmZmZmZmZmiIiIiIiIiIiId3d3VVVVZmZmVVVVZmZmZmZmZmZmd3d3ZmZmd3d3d3d3ZmZmZmZmZmZmd3d3ZmZmVVVVmZmZu7u7u7u7mZmZiIiId3d3ZmZmd3d3d3d3iIiIiIiImZmZmZmZmZmZiIiIiIiId3d3ZmZmZmZmZmZmmZmZiIiIiIiIiIiImZmZiIiId3d3iIiId3d3d3d3d3d3iIiIiIiId3d3d3d3iIiIiIiId3d3d3d3d3d3VVVVVVVVd3d3iIiIiIiId3d3REREREREVVVVVVVVREREZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREREREMzMzMzMzMzMzREREZmZmd3d3ZmZmiIiIZmZmZmZmZmZmZmZmVVVVZmZmZmZmVVVVVVVVREREREREVVVVVVVVVVVVREREREREVVVVVVVVVVVVd3d3mZmZZmZmVVVVZmZmiIiIZmZmVVVVVVVVVVVVVVVVREREREREREREZmZmZmZmVVVVVVVVZmZmVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmVVVVREREREREREREMzMzREREREREMzMzMzMzMzMzREREVVVVREREMzMzREREREREREREREREREREMzMzREREVVVVVVVVVVVVREREREREREREREREREREREREREREMzMzREREMzMzMzMzIiIiMzMzREREREREREREVVVVREREMzMzVVVVd3d3ZmZmVVVVZmZmVVVVREREREREVVVVREREREREREREREREREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVREREREREVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREVVVVMzMzMzMzMzMzIiIiMzMzIiIiIiIiERERIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzIiIiIiIiMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREREREREREREREREREREREREREREREREREMzMzVVVVVVVVZmZmZmZmREREREREREREREREREREVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREMzMzREREVVVVVVVVVVVVVVVVVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVVVVVREREVVVVVVVVVVVVVVVVREREREREREREREREVVVVd3d3d3d3ZmZmd3d3VVVVREREREREREREREREMzMzMzMzMzMzREREVVVVREREMzMzMzMzREREMzMzREREMzMzREREREREMzMzREREMzMzREREMzMzMzMzMzMzREREMzMzREREREREMzMzMzMzREREMzMzREREREREREREREREREREREREREREREREREREREREVVVVREREREREREREREREMzMzMzMzMzMzMzMzVVVVZmZmZmZmREREREREREREMzMzREREREREREREREREMzMzREREMzMzMzMzREREREREREREREREVVVVREREREREREREVVVVVVVVREREREREREREREREREREREREREREREREREREVVVVREREREREREREREREZmZmZmZmREREMzMzMzMzVVVVREREVVVVREREVVVVVVVVREREZmZmd3d3iIiImZmZVVVVMzMzREREZmZmZmZmVVVVREREREREVVVVZmZmVVVVVVVVREREVVVVREREREREVVVVZmZmVVVVVVVVZmZmREREREREREREVVVVZmZmVVVVZmZmZmZmZmZmd3d3ZmZmd3d3d3d3d3d3REREZmZmqqqq3d3d3d3d3d3d3d3dqqqqiIiIiIiIiIiImZmZiIiIiIiId3d3VVVVZmZmZmZmVVVVVVVVVVVVd3d3mZmZd3d3VVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVREREVVVVREREREREVVVVVVVViIiIqqqqd3d3VVVVVVVVREREVVVVREREiIiIqqqqiIiIVVVVVVVVmZmZzMzMzMzMu7u7qqqqmZmZiIiImZmZiIiIZmZmd3d3iIiImZmZmZmZiIiIiIiIiIiIzMzMqqqqZmZmVVVViIiIqqqqmZmZiIiIZmZmd3d3VVVVREREVVVVREREREREREREREREZmZmmZmZiIiIiIiIiIiImZmZiIiIiIiIqqqqzMzMqqqqd3d3mZmZu7u73d3d////////////////////////////////////////////7u7u//////////////////////////////////////////////////8A//8AAP////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////3d3du7u7qqqqu7u7zMzM3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u7u7u7u7u3d3d7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM3d3dzMzMzMzMzMzMzMzMzMzM3d3dzMzM3d3dzMzMzMzM3d3dzMzM3d3dzMzM3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM3d3dzMzMu7u7zMzMu7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqqqqqmZmZqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqmZmZmZmZmZmZiIiIiIiIiIiId3d3ZmZmZmZmZmZmZmZmVVVVVVVVREREREREREREREREREREREREREREREREMzMzMzMzMzMzREREMzMzREREMzMzMzMzREREREREREREREREVVVVREREREREREREREREREREVVVVVVVVVVVVREREREREREREVVVVZmZmVVVVVVVVVVVVZmZmVVVVZmZmVVVVZmZmd3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVVVVVVVVVVVVVVVVVREREREREREREREREVVVVd3d3VVVVZmZmd3d3d3d3qqqqmZmZiIiIiIiIqqqqiIiIZmZmd3d3iIiId3d3d3d3iIiIqqqqqqqqmZmZiIiImZmZd3d3d3d3d3d3d3d3d3d3d3d3VVVVZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmVVVVREREREREREREMzMzVVVVZmZmZmZmiIiIqqqqmZmZiIiIiIiImZmZzMzM3d3dzMzMzMzMzMzM3d3du7u7iIiIiIiImZmZmZmZmZmZqqqqu7u7zMzM3d3dzMzMu7u7qqqqqqqqmZmZmZmZmZmZd3d3d3d3iIiIiIiIZmZmREREZmZmd3d3d3d3qqqqqqqqmZmZiIiImZmZmZmZqqqqmZmZmZmZiIiIiIiIiIiImZmZiIiIVVVVREREVVVVREREVVVVREREZmZmd3d3VVVVREREVVVVVVVVVVVVREREREREMzMzREREREREREREREREREREVVVVREREMzMzVVVVmZmZmZmZiIiImZmZqqqqqqqqmZmZiIiId3d3d3d3ZmZmVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVZmZmd3d3iIiImZmZqqqqiIiId3d3d3d3VVVVZmZmVVVVVVVVVVVVREREVVVVREREREREVVVVREREREREZmZmmZmZmZmZiIiId3d3VVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3VVVVZmZmd3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVZmZmd3d3d3d3ZmZmd3d3d3d3d3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmd3d3VVVVVVVVd3d3mZmZqqqqqqqqmZmZiIiImZmZqqqqqqqqiIiImZmZmZmZmZmZmZmZmZmZiIiImZmZd3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmd3d3ZmZmd3d3qqqqmZmZiIiIZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmd3d3d3d3d3d3ZmZmd3d3d3d3ZmZmZmZmiIiIqqqqqqqqmZmZiIiIiIiId3d3iIiIiIiIiIiImZmZmZmZmZmZiIiIiIiId3d3ZmZmZmZmZmZmVVVVd3d3iIiIiIiImZmZmZmZd3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3VVVVVVVVd3d3mZmZmZmZd3d3ZmZmVVVVREREVVVVVVVVd3d3d3d3VVVVVVVVVVVVVVVVREREVVVVREREREREREREVVVVVVVVVVVVd3d3ZmZmd3d3ZmZmd3d3VVVVZmZmZmZmZmZmZmZmVVVVREREVVVVVVVVVVVVZmZmVVVVVVVVVVVVREREVVVVVVVVZmZmd3d3ZmZmVVVVVVVVZmZmVVVVVVVVVVVVREREREREVVVVREREZmZmZmZmVVVVZmZmZmZmVVVVVVVVREREREREZmZmREREVVVVZmZmVVVVVVVVVVVVREREVVVVREREREREREREMzMzMzMzMzMzVVVVVVVVREREREREREREREREMzMzREREMzMzREREREREREREVVVVVVVVREREREREVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVREREREREREREREREVVVVREREREREMzMzREREREREVVVVVVVVREREREREMzMzREREREREREREREREREREREREVVVVVVVVZmZmVVVVREREREREVVVVREREREREIiIiMzMzMzMzMzMzIiIiIiIiERERIiIiIiIiIiIiMzMzMzMzIiIiMzMzMzMzIiIiIiIiIiIiMzMzREREMzMzMzMzMzMzMzMzMzMzREREREREREREREREVVVVREREREREVVVVREREREREREREREREMzMzREREREREREREMzMzREREVVVVVVVVVVVVREREREREREREVVVVVVVVREREREREMzMzREREMzMzMzMzMzMzMzMzREREMzMzMzMzREREREREVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVREREREREREREMzMzREREREREMzMzMzMzREREREREVVVVVVVVVVVVVVVVREREREREVVVVREREREREVVVVVVVVVVVViIiId3d3ZmZmVVVVZmZmVVVVVVVVVVVVZmZmMzMzMzMzMzMzZmZmZmZmREREMzMzMzMzREREREREMzMzREREREREMzMzREREMzMzREREREREMzMzREREMzMzMzMzMzMzMzMzREREMzMzREREREREVVVVREREREREVVVVVVVVVVVVREREREREREREVVVVREREREREREREMzMzREREREREREREMzMzREREREREZmZmd3d3ZmZmVVVVREREVVVVREREMzMzREREMzMzMzMzMzMzREREMzMzREREREREREREREREREREREREREREVVVVREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVREREREREVVVVREREREREREREREREREREVVVVZmZmREREMzMzMzMzVVVVVVVVREREREREREREREREVVVViIiImZmZqqqqqqqqZmZmREREREREVVVVZmZmREREREREMzMzVVVVZmZmZmZmREREREREREREREREREREVVVVVVVVVVVVREREVVVVVVVVREREVVVVVVVVVVVVVVVVd3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3REREREREmZmZzMzMzMzMu7u7u7u7mZmZiIiIiIiImZmZmZmZqqqqmZmZd3d3ZmZmiIiImZmZd3d3VVVVZmZmmZmZqqqqZmZmVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmiIiId3d3ZmZmZmZmVVVVVVVVVVVVVVVVREREREREVVVVREREREREiIiIzMzMmZmZVVVVVVVVVVVVVVVVVVVVZmZmqqqqiIiIVVVVREREiIiIqqqqu7u7mZmZmZmZiIiId3d3d3d3iIiId3d3iIiImZmZiIiIiIiIiIiId3d3VVVVmZmZmZmZZmZmZmZmZmZmmZmZqqqqqqqqd3d3ZmZmZmZmVVVVVVVVREREREREMzMzVVVVVVVVZmZmd3d3d3d3iIiIiIiIiIiIiIiIiIiIu7u7u7u7iIiId3d3iIiIqqqqzMzM3d3d////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////+7u7t3d3czMzLu7u7u7u8zMzLu7u8zMzMzMzMzMzMzMzN3d3d3d3d3d3czMzMzMzN3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3d3d3e7u7t3d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3czMzN3d3czMzN3d3d3d3czMzMzMzLu7u8zMzMzMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u6qqqqqqqqqqqqqqqpmZmaqqqpmZmZmZmZmZmZmZmZmZmZmZmaqqqpmZmZmZmZmZmZmZmZmZmZmZmZmZmaqqqpmZmZmZmZmZmaqqqpmZmZmZmZmZmXd3d4iIiHd3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVURERERERERERERERDMzM0RERDMzM0RERERERDMzMzMzM0RERERERERERFVVVURERERERERERFVVVURERERERERERERERERERERERERERDMzM0RERERERERERERERFVVVURERERERERERERERERERERERERERFVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERDMzM0RERERERFVVVVVVVVVVVWZmZmZmZoiIiKqqqpmZmYiIiIiIiIiIiGZmZlVVVXd3d3d3d4iIiHd3d3d3d5mZmaqqqoiIiJmZmYiIiHd3d3d3d2ZmZnd3d4iIiHd3d1VVVWZmZmZmZnd3d3d3d2ZmZmZmZmZmZmZmZmZmZlVVVWZmZkRERERERERERERERGZmZmZmZlVVVYiIiKqqqoiIiIiIiIiIiKqqqszMzN3d3bu7u7u7u8zMzMzMzIiIiHd3d5mZmZmZmYiIiIiIiKqqqpmZmczMzN3d3czMzKqqqqqqqqqqqpmZmYiIiIiIiHd3d3d3d4iIiHd3d0RERFVVVWZmZnd3d4iIiJmZmaqqqpmZmYiIiJmZmaqqqqqqqpmZmYiIiIiIiIiIiIiIiIiIiGZmZlVVVWZmZmZmZmZmZmZmZlVVVVVVVXd3d2ZmZlVVVURERGZmZmZmZkRERFVVVURERERERERERFVVVVVVVVVVVVVVVVVVVVVVVURERIiIiKqqqpmZmZmZmZmZmYiIiHd3d2ZmZmZmZnd3d1VVVURERFVVVWZmZmZmZlVVVVVVVWZmZlVVVURERGZmZoiIiJmZmZmZmZmZmWZmZnd3d2ZmZlVVVURERFVVVVVVVVVVVURERERERERERERERFVVVURERERERGZmZoiIiIiIiHd3d2ZmZlVVVVVVVWZmZlVVVVVVVWZmZmZmZmZmZmZmZlVVVWZmZnd3d4iIiGZmZlVVVWZmZmZmZnd3d3d3d3d3d2ZmZmZmZnd3d3d3d3d3d4iIiGZmZnd3d3d3d2ZmZlVVVVVVVVVVVVVVVXd3d3d3d3d3d2ZmZnd3d3d3d3d3d3d3d2ZmZnd3d2ZmZlVVVVVVVWZmZmZmZkRERFVVVYiIiIiIiJmZmaqqqpmZmZmZmYiIiJmZmYiIiJmZmZmZmYiIiIiIiIiIiIiIiHd3d4iIiIiIiHd3d4iIiHd3d3d3d2ZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZnd3d2ZmZoiIiKqqqqqqqoiIiHd3d2ZmZmZmZnd3d3d3d2ZmZnd3d3d3d2ZmZmZmZnd3d3d3d2ZmZoiIiIiIiHd3d2ZmZoiIiKqqqru7u6qqqoiIiIiIiIiIiIiIiIiIiIiIiJmZmZmZmYiIiJmZmYiIiHd3d2ZmZnd3d1VVVVVVVWZmZoiIiJmZmaqqqoiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiHd3d2ZmZnd3d2ZmZmZmZlVVVWZmZoiIiJmZmXd3d2ZmZkRERFVVVXd3d2ZmZnd3d2ZmZlVVVVVVVVVVVVVVVURERERERERERFVVVVVVVVVVVVVVVWZmZmZmZnd3d3d3d3d3d3d3d1VVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVVVVVVVVVURERFVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVURERERERERERFVVVVVVVWZmZmZmZlVVVWZmZmZmZlVVVURERERERERERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERDMzMzMzMzMzM0RERFVVVURERERERERERDMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERFVVVVVVVURERERERERERDMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVTMzM0RERDMzM0RERERERERERERERFVVVWZmZmZmZmZmZlVVVVVVVURERERERERERFVVVVVVVVVVVURERDMzM0RERERERFVVVVVVVURERDMzM0RERDMzM0RERDMzM0RERERERERERERERFVVVWZmZkRERERERERERERERDMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIjMzMyIiIiIiIjMzMzMzMzMzMyIiIiIiIjMzM0RERERERFVVVVVVVURERFVVVURERDMzM0RERFVVVURERERERERERDMzM0RERDMzM0RERERERDMzM0RERERERERERERERFVVVVVVVWZmZkRERERERERERDMzMzMzMzMzMzMzM0RERERERDMzMzMzM0RERDMzM1VVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERDMzMzMzM0RERDMzMzMzM0RERERERFVVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVURERGZmZoiIiKqqqmZmZlVVVVVVVVVVVWZmZnd3d1VVVTMzMzMzM0RERHd3d2ZmZkRERDMzMzMzMzMzM0RERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERFVVVVVVVVVVVVVVVURERERERERERFVVVVVVVVVVVURERERERDMzM0RERERERERERERERERERERERGZmZmZmZmZmZlVVVURERERERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERERERERERERERERERFVVVURERERERFVVVURERFVVVVVVVVVVVVVVVURERERERDMzM0RERDMzM0RERERERERERFVVVURERFVVVURERDMzMzMzM0RERERERERERDMzM0RERDMzM1VVVYiIiIiIiLu7u5mZmVVVVURERERERGZmZnd3d0RERERERDMzM0RERFVVVVVVVURERERERERERERERERERFVVVURERERERERERFVVVVVVVVVVVVVVVWZmZlVVVVVVVWZmZnd3d2ZmZnd3d2ZmZmZmZnd3d4iIiERERERERIiIiLu7u7u7u5mZmaqqqpmZmYiIiHd3d4iIiJmZmaqqqqqqqoiIiHd3d4iIiKqqqoiIiGZmZlVVVXd3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVURERFVVVWZmZqqqqszMzIiIiERERERERERERFVVVVVVVXd3d5mZmYiIiFVVVVVVVYiIiLu7u6qqqoiIiJmZmYiIiHd3d2ZmZnd3d3d3d4iIiIiIiHd3d3d3d3d3d3d3d1VVVWZmZlVVVVVVVVVVVWZmZoiIiJmZmbu7u4iIiGZmZlVVVURERERERERERERERERERERERFVVVWZmZlVVVWZmZnd3d2ZmZoiIiIiIiHd3d5mZmbu7u4iIiGZmZnd3d3d3d5mZmczMzN3d3f///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////u7u7d3d3d3d3MzMzMzMzMzMzMzMzd3d3MzMzd3d3MzMzMzMzMzMzd3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3d3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzd3d3MzMzd3d3MzMy7u7vMzMzMzMzMzMy7u7vMzMy7u7u7u7u7u7uqqqqqqqqZmZmZmZmZmZmIiIiIiIiZmZmZmZmZmZmZmZmZmZmqqqqZmZmZmZmIiIiIiIiZmZmZmZmZmZmZmZmZmZmqqqqZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmIiIiIiIiIiIh3d3dmZmZ3d3dmZmZVVVVERERVVVVEREREREREREQzMzMzMzNEREREREREREREREREREREREREREREREREREQzMzNEREREREQzMzNERERERERERERERERVVVVmZmZVVVVVVVVVVVUzMzMzMzNVVVVEREREREQzMzMzMzNEREQzMzNERERERERERERVVVVVVVVERERERERERERVVVVmZmZERERERERERERERERVVVVERERERERERERVVVVmZmaIiIiZmZl3d3dmZmZmZmZmZmZERERVVVV3d3eIiIiIiIh3d3eIiIiZmZmIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZVVVVVVVV3d3eIiIh3d3dmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVWIiIiZmZmIiIiIiIiIiIiqqqrd3d3d3d3MzMyqqqqqqqq7u7uZmZmIiIiZmZmZmZl3d3d3d3d3d3d3d3e7u7vMzMzMzMy7u7u7u7uZmZmZmZmIiIiIiIh3d3eIiIiIiIh3d3d3d3d3d3eZmZmIiIh3d3eIiIiqqqqZmZmIiIiIiIiZmZmIiIiZmZmIiIiIiIiIiIiIiIiIiIh3d3dmZmZ3d3eIiIh3d3d3d3dVVVVERERmZmZ3d3dmZmZERERmZmZmZmZERERERERVVVVmZmZmZmZmZmZVVVVERERmZmZmZmZmZmZmZmZ3d3eIiIiZmZmZmZmZmZmIiIhmZmZVVVVmZmZVVVVVVVVVVVVmZmZVVVVmZmZVVVVERERVVVVVVVVmZmZmZmZmZmaIiIiIiIh3d3d3d3dmZmZmZmZVVVVVVVVmZmZmZmZVVVVVVVVVVVVERERERERVVVVVVVVERERERER3d3eIiIhmZmZmZmZmZmZVVVVmZmZVVVVVVVVVVVV3d3dmZmZmZmZmZmZ3d3dmZmaIiIh3d3dVVVVVVVVVVVV3d3d3d3d3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dVVVVERERVVVWIiIiIiIiIiIiIiIiIiIiIiIhmZmZ3d3d3d3d3d3dmZmZmZmZVVVVmZmZVVVVERERERESIiIiZmZmZmZmqqqqZmZmZmZmIiIiIiIiIiIiZmZmIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3eIiIiIiIh3d3dmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3eZmZmZmZl3d3d3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3dmZmZ3d3d3d3dmZmaIiIi7u7u7u7uqqqqZmZmIiIiIiIh3d3d3d3eZmZmIiIiZmZmIiIiIiIiIiIiIiIiIiIh3d3dVVVVVVVVmZmaIiIiZmZmZmZmqqqqIiIh3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIh3d3d3d3d3d3dmZmZmZmZVVVVVVVVmZmaIiIiZmZl3d3dVVVVERERmZmZ3d3dmZmZVVVVERERVVVVERERVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVV3d3d3d3eIiIhmZmZVVVVVVVVVVVVVVVVERERERERVVVVmZmZmZmZ3d3dVVVVERERERERERERVVVVVVVVVVVVVVVVVVVV3d3dmZmZmZmZmZmZVVVVERERERERERERERERVVVVmZmZmZmZmZmZmZmZmZmZVVVVEREREREREREQzMzNERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVEREREREQzMzMzMzMzMzNERERVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVVVVVEREQzMzNEREREREREREREREQzMzMzMzNERERERERVVVVVVVVVVVVEREQzMzNERERERERVVVVERERVVVVVVVV3d3dmZmZmZmZVVVVVVVVERERERERERERVVVVVVVVVVVVERERVVVVVVVVVVVVEREREREQzMzNEREREREREREQzMzNERERERERERERERERVVVVVVVVVVVVVVVVVVVUzMzMiIiIiIiIiIiIzMzMzMzMiIiIREREiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIzMzMzMzMzMzMiIiIiIiIzMzNERERVVVVERERVVVVVVVVEREREREQzMzNEREREREREREREREREREREREQzMzNERERERERERERERERVVVVERERERERERERERERmZmZVVVVVVVVEREREREREREREREQzMzNEREQzMzMzMzNEREQzMzMzMzNERERERERERERERERVVVVERERERERVVVVVVVVVVVUzMzNEREREREREREREREQzMzMzMzMzMzMzMzNERERERERERERVVVVVVVVVVVVVVVVERERVVVVVVVVERERERER3d3eqqqqqqqp3d3dVVVVVVVVVVVVmZmZ3d3dVVVUzMzMzMzMzMzNmZmZmZmYzMzMzMzMzMzMzMzMzMzMiIiIzMzNEREQzMzNEREREREQzMzNEREQzMzMzMzNEREQzMzMzMzMzMzNERERERERERERERERVVVVERERVVVVVVVVERERVVVVERERVVVVVVVVEREREREREREQzMzNEREQzMzMzMzNERERERERERERVVVVEREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERERERERERERERERERERERERERERERERERERERVVVVVVVVVVVUzMzNEREQzMzMzMzMzMzMzMzNERERVVVVERERERERVVVVmZmZEREQzMzNEREREREREREREREQzMzNERERVVVVmZmZ3d3e7u7uZmZlVVVVERERERER3d3eZmZlVVVVEREQzMzNERERVVVVEREQzMzMzMzMzMzNERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3dmZmZmZmaIiIhVVVUzMzNmZma7u7uqqqqqqqqZmZmZmZmIiIh3d3eIiIiIiIiZmZmIiIiZmZmIiIiIiIiZmZmqqqqqqqp3d3dERERmZmZ3d3dVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmaZmZnMzMy7u7t3d3dERERVVVVERERERERERER3d3eqqqqqqqpVVVVERER3d3e7u7uqqqqZmZmqqqqZmZl3d3dmZmZmZmZmZmaIiIiIiIh3d3eZmZmIiIiIiIh3d3dmZmZVVVVVVVVmZmZmZmZmZmaqqqrMzMzMzMyIiIhVVVVVVVVVVVVVVVVERERERERERERVVVVVVVVmZmZmZmZmZmZmZmZ3d3eIiIh3d3eIiIiqqqqZmZlmZmZVVVVmZmaIiIiZmZm7u7vd3d3u7u7////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzM3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzMzMzMzMzM3d3dzMzMzMzMzMzMzMzMu7u7u7u7zMzMzMzMu7u7u7u7qqqqqqqqmZmZqqqqmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZiIiImZmZmZmZmZmZmZmZqqqqmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZiIiImZmZiIiIiIiIiIiIiIiId3d3ZmZmZmZmZmZmVVVVREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREMzMzREREREREVVVVZmZmZmZmVVVVVVVVZmZmVVVVMzMzVVVVZmZmVVVVREREREREREREREREMzMzREREREREREREVVVVVVVVREREVVVVVVVVZmZmZmZmREREREREREREVVVVZmZmVVVVREREREREREREVVVVVVVVZmZmZmZmVVVVVVVVVVVVREREREREZmZmiIiId3d3iIiImZmZiIiId3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmVVVVREREVVVVd3d3d3d3ZmZmZmZmZmZmVVVVREREREREVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3ZmZmd3d3ZmZmiIiImZmZmZmZu7u77u7u3d3dzMzMu7u7qqqqqqqqqqqqmZmZmZmZiIiId3d3d3d3iIiIiIiIqqqqu7u73d3du7u7qqqqmZmZmZmZmZmZiIiId3d3iIiImZmZiIiImZmZqqqqqqqqmZmZiIiIiIiImZmZqqqqiIiId3d3d3d3iIiId3d3iIiIiIiId3d3d3d3iIiId3d3d3d3iIiId3d3d3d3d3d3ZmZmVVVVVVVVd3d3d3d3ZmZmZmZmVVVVREREREREZmZmd3d3d3d3d3d3ZmZmVVVVVVVVVVVVVVVVd3d3ZmZmd3d3iIiIiIiIiIiIiIiId3d3d3d3ZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3ZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVVVVVREREVVVVVVVVd3d3d3d3ZmZmd3d3ZmZmZmZmd3d3iIiIVVVVVVVVZmZmd3d3ZmZmVVVVVVVVd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIZmZmVVVVREREZmZmmZmZiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3ZmZmZmZmVVVVd3d3ZmZmVVVVVVVVd3d3mZmZqqqqqqqqqqqqmZmZmZmZd3d3d3d3mZmZmZmZiIiImZmZiIiIiIiId3d3ZmZmd3d3d3d3iIiId3d3ZmZmVVVVZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiIiIiId3d3d3d3ZmZmZmZmd3d3d3d3mZmZiIiId3d3iIiIZmZmd3d3ZmZmd3d3iIiIiIiId3d3d3d3d3d3ZmZmd3d3d3d3ZmZmZmZmZmZmZmZmiIiIu7u7u7u7u7u7iIiIiIiIiIiIiIiIiIiImZmZiIiId3d3iIiId3d3iIiImZmZiIiIVVVVVVVVREREVVVVmZmZmZmZqqqqmZmZiIiId3d3d3d3d3d3d3d3iIiImZmZiIiIiIiIiIiId3d3d3d3iIiIZmZmVVVVVVVVZmZmd3d3iIiIiIiId3d3ZmZmVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVREREREREVVVVVVVVZmZmZmZmREREREREVVVVVVVVZmZmZmZmiIiId3d3VVVVVVVVVVVVVVVVREREREREREREVVVVd3d3d3d3ZmZmZmZmREREMzMzREREVVVVVVVVREREREREVVVVZmZmZmZmVVVVZmZmVVVVREREMzMzREREVVVVVVVVZmZmZmZmZmZmZmZmVVVVVVVVREREREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVMzMzREREMzMzREREMzMzREREVVVVVVVVREREREREMzMzMzMzIiIiMzMzREREMzMzMzMzMzMzMzMzREREVVVVVVVVREREVVVVREREREREREREREREREREREREREREVVVVVVVVVVVVREREREREREREREREVVVVZmZmVVVVREREVVVVZmZmVVVVVVVVVVVVVVVVREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREMzMzREREREREMzMzREREVVVVREREREREVVVVREREVVVVREREMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiERERIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzIiIiIiIiMzMzIiIiMzMzREREREREREREVVVVREREREREMzMzMzMzREREREREREREREREREREMzMzMzMzREREREREREREVVVVVVVVVVVVREREREREVVVVZmZmVVVVVVVVVVVVREREREREMzMzREREMzMzREREREREMzMzMzMzMzMzREREREREREREREREZmZmREREREREREREVVVVREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVREREVVVVmZmZzMzMqqqqZmZmVVVVd3d3d3d3ZmZmd3d3VVVVMzMzIiIiMzMzVVVVVVVVMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiMzMzREREMzMzREREMzMzMzMzMzMzREREMzMzREREREREREREREREREREREREVVVVVVVVREREREREREREVVVVREREVVVVVVVVREREREREREREREREREREREREREREREREREREMzMzREREREREMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREVVVVREREREREREREREREREREMzMzREREMzMzREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVREREREREZmZmVVVVMzMzREREREREREREREREMzMzMzMzVVVVZmZmiIiIqqqqqqqqVVVVVVVVVVVVd3d3iIiIVVVVREREMzMzREREREREMzMzREREMzMzREREREREREREREREMzMzREREVVVVVVVVREREREREVVVVVVVVVVVVVVVVZmZmVVVVZmZmiIiId3d3ZmZmZmZmd3d3VVVVMzMzVVVVmZmZmZmZiIiImZmZmZmZd3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3iIiIiIiIqqqqzMzMqqqqZmZmZmZmd3d3VVVVREREREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmu7u77u7uqqqqZmZmREREREREREREVVVVVVVViIiIzMzMmZmZREREREREmZmZu7u7qqqqu7u7qqqqiIiId3d3ZmZmVVVVZmZmiIiId3d3d3d3mZmZqqqqiIiImZmZd3d3VVVVVVVVZmZmVVVVZmZmmZmZzMzM3d3dzMzMmZmZZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmd3d3iIiIiIiId3d3d3d3mZmZu7u7d3d3VVVVVVVVZmZmd3d3mZmZu7u77u7u////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////+7u7u7u7t3d3d3d3d3d3d3d3d3d3e7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqqqqqqqqqqqqqqqqqqqqqru7u6qqqqqqqqqqqqqqqpmZmZmZmZmZmZmZmZmZmYiIiIiIiIiIiJmZmZmZmZmZmZmZmYiIiJmZmZmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d4iIiHd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZlVVVVVVVURERDMzMzMzMzMzMzMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVURERERERFVVVURERDMzM0RERFVVVWZmZmZmZlVVVVVVVTMzMzMzM0RERGZmZmZmZkRERFVVVVVVVVVVVURERERERFVVVURERERERFVVVWZmZnd3d2ZmZkRERERERDMzM0RERDMzM0RERERERERERERERFVVVURERERERFVVVVVVVWZmZnd3d4iIiIiIiHd3d1VVVWZmZnd3d2ZmZmZmZlVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZlVVVWZmZlVVVURERFVVVVVVVVVVVURERFVVVYiIiJmZmbu7u8zMzIiIiGZmZnd3d5mZmbu7u6qqqru7u93d3czMzMzMzMzMzLu7u7u7u7u7u5mZmYiIiIiIiJmZmZmZmaqqqru7u8zMzKqqqru7u8zMzLu7u5mZmZmZmaqqqoiIiHd3d4iIiJmZmaqqqru7u6qqqpmZmYiIiIiIiJmZmZmZmZmZmZmZmYiIiIiIiIiIiGZmZnd3d3d3d2ZmZoiIiIiIiGZmZnd3d2ZmZmZmZlVVVVVVVWZmZmZmZlVVVWZmZoiIiJmZmWZmZkRERERERERERHd3d4iIiIiIiHd3d2ZmZmZmZmZmZlVVVURERFVVVURERFVVVWZmZmZmZnd3d4iIiJmZmYiIiGZmZnd3d2ZmZlVVVWZmZmZmZmZmZlVVVWZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZlVVVWZmZmZmZlVVVWZmZnd3d1VVVWZmZmZmZlVVVWZmZmZmZlVVVURERFVVVVVVVURERFVVVURERFVVVWZmZnd3d1VVVURERERERFVVVWZmZnd3d2ZmZnd3d3d3d3d3d2ZmZnd3d3d3d2ZmZlVVVXd3d3d3d1VVVVVVVWZmZnd3d3d3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d3d3d0RERERERFVVVXd3d4iIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d4iIiHd3d2ZmZlVVVWZmZoiIiGZmZlVVVXd3d5mZmaqqqqqqqoiIiIiIiJmZmYiIiJmZmYiIiJmZmZmZmaqqqoiIiHd3d3d3d2ZmZoiIiJmZmYiIiHd3d2ZmZnd3d2ZmZnd3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d2ZmZnd3d4iIiIiIiKqqqpmZmYiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d4iIiGZmZlVVVXd3d3d3d2ZmZpmZmaqqqszMzMzMzJmZmYiIiIiIiIiIiJmZmYiIiHd3d3d3d3d3d4iIiJmZmZmZmYiIiFVVVVVVVURERFVVVYiIiJmZmZmZmZmZmYiIiHd3d3d3d3d3d3d3d3d3d4iIiHd3d4iIiHd3d4iIiGZmZnd3d2ZmZmZmZmZmZmZmZnd3d3d3d4iIiHd3d2ZmZmZmZmZmZlVVVVVVVURERFVVVURERFVVVVVVVURERFVVVXd3d3d3d1VVVURERERERERERERERFVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVURERFVVVVVVVWZmZmZmZmZmZlVVVWZmZlVVVURERDMzM0RERERERERERFVVVURERERERFVVVVVVVURERERERFVVVURERDMzM1VVVVVVVWZmZnd3d2ZmZmZmZmZmZlVVVURERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVURERERERDMzM0RERERERERERFVVVVVVVVVVVVVVVURERERERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIkRERERERERERFVVVURERFVVVVVVVTMzM0RERERERFVVVVVVVVVVVVVVVURERERERDMzM0RERGZmZlVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVURERERERDMzM0RERERERERERFVVVVVVVVVVVURERFVVVURERERERDMzM0RERDMzM0RERDMzM0RERFVVVURERERERERERERERERERERERERERERERDMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERERERERERERERFVVVURERERERDMzMzMzMzMzM0RERERERERERERERERERDMzMzMzM0RERERERERERERERERERERERFVVVWZmZmZmZmZmZlVVVVVVVURERERERERERERERERERERERDMzM0RERDMzMzMzMzMzMzMzMzMzM0RERFVVVURERERERERERERERERERERERERERERERERERERERERERDMzMzMzM0RERFVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVURERERERFVVVaqqqt3d3ZmZmVVVVVVVVYiIiIiIiGZmZlVVVURERDMzMzMzMzMzM3d3d3d3d0RERCIiIjMzMyIiIiIiIiIiIhERESIiIjMzMzMzM0RERDMzM0RERDMzMzMzMzMzM0RERERERERERERERERERERERERERERERERERERERERERERERERERFVVVVVVVWZmZlVVVURERERERERERERERERERFVVVURERERERERERDMzMzMzMyIiIhERETMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM1VVVURERERERERERERERFVVVURERDMzM0RERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM1VVVWZmZlVVVTMzM0RERFVVVURERDMzM0RERDMzMzMzM0RERERERFVVVYiIiJmZmbu7u7u7u2ZmZkRERERERFVVVXd3d2ZmZkRERERERERERERERERERERERERERERERERERDMzMzMzM0RERERERFVVVURERERERERERFVVVVVVVWZmZlVVVVVVVWZmZnd3d5mZmXd3d2ZmZmZmZnd3d2ZmZjMzMzMzM2ZmZoiIiHd3d4iIiIiIiHd3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZnd3d4iIiJmZmczMzN3d3Xd3d1VVVYiIiHd3d0RERGZmZnd3d1VVVVVVVVVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVURERERERERERERERERERJmZmaqqqnd3d0RERERERFVVVVVVVVVVVVVVVZmZmczMzHd3d0RERERERIiIiJmZmbu7u8zMzIiIiHd3d3d3d2ZmZnd3d3d3d3d3d2ZmZmZmZoiIiLu7u6qqqoiIiHd3d3d3d1VVVURERERERFVVVVVVVYiIiMzMzO7u7u7u7szMzIiIiFVVVURERERERERERGZmZlVVVVVVVURERHd3d4iIiHd3d4iIiHd3d3d3d4iIiKqqqpmZmXd3d0RERERERERERFVVVYiIiLu7u93d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7u7u7d3d3u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3d3d3u7u7d3d3u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3MzMzMzMzMzMy7u7u7u7u7u7u7u7uqqqq7u7uqqqqqqqqqqqqZmZmqqqqZmZmZmZmqqqqZmZmqqqqqqqqqqqqZmZmZmZmZmZmZmZmZmZmZmZmIiIiZmZmIiIiZmZmZmZmIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3eIiIh3d3eIiIiIiIh3d3d3d3d3d3eIiIh3d3d3d3dmZmZ3d3dmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVEREREREREREQzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzNERERERERVVVVVVVVEREQzMzNERERVVVVVVVVERERVVVVVVVVVVVVVVVVEREREREREREQzMzNERERERERVVVVmZmZERERERERVVVVmZmZVVVVVVVVVVVVEREQzMzNERERERERERERERERVVVVVVVVmZmZ3d3dmZmZmZmZmZmZmZmZVVVVmZmZ3d3dmZmZVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERESIiIiZmZnMzMzd3d2ZmZl3d3eZmZm7u7u7u7uqqqq7u7vd3d3MzMzd3d3MzMzMzMy7u7uqqqqZmZmIiIiZmZm7u7u7u7uqqqrMzMy7u7u7u7uqqqq7u7u7u7uZmZmqqqqqqqqZmZmZmZmZmZmZmZmqqqqqqqqZmZmZmZmIiIiIiIiIiIh3d3eIiIiZmZmZmZmIiIh3d3dmZmZ3d3dmZmZmZmaIiIiIiIh3d3d3d3dmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZ3d3eIiIh3d3dEREQzMzNVVVWIiIiIiIiIiIhmZmZmZmZVVVVVVVVmZmZVVVVVVVVERERERERmZmZmZmZVVVVmZmaIiIh3d3dmZmZmZmZVVVVmZmZmZmZmZmZVVVVmZmZVVVVmZmZ3d3dmZmZmZmZVVVVmZmZVVVVERERVVVVmZmZmZmZmZmZVVVVmZmZmZmZmZmZ3d3eIiIh3d3dVVVVERERERERERERVVVVVVVVERERERER3d3dmZmZmZmZVVVVVVVVVVVVmZmZ3d3d3d3d3d3dmZmZ3d3dmZmZ3d3d3d3dVVVVVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3eIiIiIiIh3d3d3d3d3d3d3d3dVVVVERERmZmaIiIiIiIiIiIiIiIiIiIiIiIiZmZmIiIh3d3eIiIiIiIhmZmZVVVVVVVWIiIhVVVVVVVV3d3eZmZmqqqqZmZmIiIiIiIiZmZmZmZmZmZmZmZmIiIiZmZmqqqqZmZmIiIiIiIh3d3eZmZmZmZmIiIh3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIi7u7uqqqqZmZmIiIh3d3d3d3d3d3dmZmZmZmZmZmZ3d3d3d3dmZmZmZmaIiIh3d3dmZmZ3d3d3d3dmZmZmZmaqqqq7u7u7u7uZmZmIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZmIiIiIiIh3d3dmZmZmZmZmZmZmZmZ3d3eZmZmZmZmIiIiIiIh3d3eIiIhmZmZVVVV3d3d3d3d3d3d3d3d3d3eIiIh3d3dmZmZmZmZmZmZmZmZVVVVmZmZmZmZ3d3d3d3dmZmZVVVV3d3d3d3dVVVVVVVVERERERERVVVVERERVVVVmZmZ3d3dmZmZmZmZERERERERERERERERVVVVERERVVVVVVVVmZmZERERVVVVERERERERERERmZmZ3d3d3d3dVVVVmZmZmZmZVVVVEREQzMzMzMzNVVVVVVVVVVVVERERVVVVVVVVVVVVEREREREREREREREQzMzNERERVVVV3d3dmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERVVVVVVVVVVVVEREQzMzNERERVVVVVVVVVVVVVVVVVVVVVVVVEREREREREREREREREREQzMzMzMzMiIiIzMzNEREQzMzMzMzMzMzNERERERERERERERERVVVVERERERERERERERERERERVVVVVVVVEREREREREREQzMzNERERERERVVVVERERERERERERERERVVVVVVVVEREREREREREQzMzMzMzMzMzNERERVVVVVVVVVVVVERERVVVVEREREREREREQzMzNEREREREQzMzNERERERERVVVVEREQzMzNEREREREREREREREREREQzMzMzMzMiIiIiIiIiIiIzMzMiIiIREREiIiIiIiIzMzMiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzNERERERERVVVVERERVVVVEREQzMzNEREREREREREREREREREREREQzMzNEREQzMzMzMzNEREREREQzMzNEREQzMzNERERVVVVmZmZVVVVmZmZmZmZEREREREREREREREQzMzNEREQzMzNEREQzMzNEREQzMzMzMzNEREQzMzNERERERERERERERERERERERERVVVVEREQzMzNEREQzMzMzMzMzMzMzMzNERERERERERERVVVVmZmZVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVWZmZm7u7uIiIhVVVVERER3d3d3d3dmZmZVVVVEREQzMzMzMzMzMzN3d3d3d3dEREQzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiJEREQzMzNEREQzMzNEREQzMzNEREQzMzNERERERERERERERERERERERERERERERERERERERERERERERERVVVVVVVVVVVVEREREREREREREREREREREREREREREREQzMzMzMzMzMzMiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMiIiIzMzMzMzNERERERERERERERERVVVVERERERERERERVVVVEREREREREREQzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzNERERERERERESIiIhVVVVERERERERERERVVVVEREQzMzMzMzNEREQzMzNERERVVVV3d3eIiIiqqqqqqqpVVVVERERERERVVVVmZmZmZmZERERERERVVVVVVVVVVVUzMzMzMzMzMzMzMzMzMzNEREQzMzNVVVVVVVVVVVVERERERERmZmZVVVVmZmZVVVVVVVVmZmZmZmaIiIh3d3dmZmZ3d3d3d3d3d3dEREQiIiJVVVV3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZ3d3eIiIiqqqrMzMx3d3dVVVV3d3d3d3dVVVVmZmZ3d3dVVVVVVVVERERERERERERERERERERERERVVVVmZmZVVVVVVVVmZmZVVVVVVVVERERERERERERERERERERERERVVVVmZmZmZmZVVVVERERVVVVERERVVVVVVVVmZmaqqqqqqqpmZmZERERERESIiIiqqqq7u7uqqqqIiIh3d3d3d3d3d3eIiIh3d3dmZmZmZmZmZmZ3d3eqqqqqqqp3d3d3d3eIiIiIiIhVVVVmZmZVVVVVVVVmZmaIiIjMzMzu7u7d3d2qqqp3d3dVVVVERERERERVVVVERERERERVVVWZmZmIiIh3d3d3d3d3d3d3d3d3d3eZmZmqqqp3d3dVVVVERERERERERERmZmaZmZm7u7vMzMzu7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMu7u7u7u7qqqqqqqqqqqqu7u7u7u7u7u7u7u7qqqqqqqqu7u7u7u7u7u7zMzMzMzMzMzM3d3dzMzMzMzM3d3dzMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3dzMzM3d3d3d3d3d3dzMzM3d3dzMzM3d3dzMzM3d3dzMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7qqqqu7u7qqqqqqqqqqqqqqqqmZmZmZmZmZmZmZmZmZmZmZmZmZmZqqqqmZmZqqqqmZmZqqqqmZmZqqqqmZmZmZmZiIiIiIiIiIiIiIiIiIiId3d3iIiIiIiId3d3d3d3d3d3iIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3ZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmREREVVVVVVVVREREREREREREVVVVVVVVREREVVVVMzMzREREMzMzREREMzMzMzMzREREMzMzMzMzMzMzREREREREREREMzMzMzMzREREVVVVVVVVREREREREVVVVVVVVREREREREREREREREREREREREREREVVVVVVVVREREVVVVZmZmZmZmVVVVZmZmVVVVMzMzMzMzMzMzMzMzREREREREZmZmd3d3d3d3VVVVZmZmVVVVVVVVVVVVZmZmZmZmd3d3ZmZmVVVVVVVVVVVVZmZmVVVVZmZmREREREREVVVVVVVVVVVVVVVVREREREREREREREREiIiImZmZzMzM7u7uzMzMd3d3mZmZzMzMu7u7qqqqu7u7zMzM3d3dzMzMzMzMzMzMzMzMqqqqqqqqmZmZu7u7zMzMqqqqqqqqu7u7zMzMqqqqmZmZu7u7u7u7qqqqqqqqqqqqmZmZqqqqmZmZmZmZiIiImZmZiIiIiIiIiIiIiIiIiIiId3d3d3d3iIiImZmZiIiIiIiId3d3d3d3VVVVd3d3mZmZmZmZZmZmd3d3iIiIZmZmd3d3ZmZmd3d3d3d3d3d3d3d3ZmZmd3d3d3d3ZmZmVVVVZmZmd3d3mZmZd3d3d3d3VVVVREREVVVVZmZmZmZmZmZmVVVVVVVVVVVVZmZmREREVVVVd3d3ZmZmiIiId3d3d3d3VVVVZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVd3d3iIiIREREREREZmZmVVVVZmZmVVVVVVVVVVVVVVVVZmZmmZmZiIiIZmZmVVVVVVVVVVVVREREREREVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmREREVVVVZmZmd3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3iIiId3d3ZmZmREREVVVVmZmZmZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIZmZmZmZmZmZmVVVVd3d3VVVVVVVViIiIqqqqu7u7mZmZiIiIqqqqqqqqmZmZmZmZmZmZmZmZmZmZiIiImZmZmZmZmZmZiIiIiIiImZmZiIiId3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3ZmZmd3d3d3d3iIiIqqqqu7u7mZmZd3d3iIiId3d3d3d3ZmZmZmZmZmZmd3d3ZmZmd3d3d3d3iIiIZmZmVVVVZmZmd3d3VVVVVVVViIiIzMzMu7u7mZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZmZmZiIiId3d3ZmZmd3d3d3d3iIiIiIiId3d3iIiImZmZmZmZiIiId3d3iIiIZmZmVVVVd3d3ZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmREREREREREREREREREREREREREREVVVVREREREREVVVVREREMzMzREREd3d3d3d3iIiId3d3ZmZmd3d3ZmZmREREREREREREREREREREREREVVVVVVVVREREREREMzMzREREREREMzMzREREVVVVVVVVd3d3d3d3ZmZmVVVVZmZmVVVVREREVVVVREREREREREREREREREREREREREREREREREREVVVVREREREREVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzREREMzMzREREVVVVVVVVREREVVVVVVVVREREREREVVVVREREREREREREREREREREREREVVVVREREREREMzMzREREVVVVVVVVREREREREREREREREMzMzREREVVVVVVVVVVVVVVVVVVVVREREMzMzREREMzMzREREREREMzMzREREREREREREVVVVREREREREMzMzMzMzREREREREMzMzMzMzIiIiMzMzIiIiMzMzIiIiIiIiERERIiIiIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzREREREREVVVVREREVVVVREREREREREREREREREREREREVVVVREREREREREREREREMzMzMzMzREREREREMzMzMzMzMzMzMzMzZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREREREREREREREREREMzMzREREMzMzREREREREREREREREREREVVVVREREREREREREMzMzREREREREMzMzREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVZmZmd3d3iIiId3d3VVVVVVVVVVVVZmZmZmZmZmZmREREMzMzMzMzMzMzVVVVd3d3VVVVMzMzMzMzIiIiIiIiIiIiMzMzIiIiIiIiMzMzMzMzMzMzREREMzMzMzMzMzMzREREREREREREREREREREREREREREREREREREVVVVREREREREREREVVVVREREREREVVVVREREREREREREREREVVVVREREMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiREREREREVVVVREREREREREREMzMzREREVVVVVVVVVVVVREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREZmZmVVVVREREMzMzREREVVVVREREREREMzMzMzMzREREREREZmZmZmZmd3d3mZmZmZmZVVVVREREREREREREZmZmZmZmREREREREVVVVVVVVREREMzMzMzMzMzMzMzMzMzMzREREREREVVVVVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVZmZmd3d3d3d3d3d3d3d3iIiId3d3d3d3ZmZmIiIiREREd3d3ZmZmd3d3ZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmZmZmd3d3mZmZd3d3VVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVREREVVVVMzMzREREVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVREREVVVVREREREREREREREREREREVVVVVVVVd3d3ZmZmREREVVVVVVVVVVVVZmZmmZmZiIiIVVVVMzMzVVVVqqqqu7u7u7u7mZmZd3d3d3d3d3d3d3d3d3d3d3d3ZmZmVVVVZmZmd3d3mZmZzMzMmZmZd3d3ZmZmZmZmd3d3d3d3ZmZmZmZmZmZmiIiIiIiIqqqqzMzM3d3du7u7iIiIVVVVREREREREREREVVVVd3d3iIiIiIiId3d3ZmZmd3d3ZmZmZmZmiIiImZmZmZmZVVVVREREREREREREREREZmZmmZmZzMzMzMzM7u7u////////////////7u7u////////7u7u////////7u7u////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////93d3d3d3czMzN3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzLu7u7u7u6qqqqqqqqqqqru7u7u7u7u7u6qqqpmZmZmZmaqqqqqqqqqqqru7u8zMzLu7u7u7u7u7u7u7u6qqqru7u6qqqqqqqqqqqqqqqqqqqru7u7u7u7u7u7u7u8zMzMzMzMzMzLu7u7u7u7u7u8zMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqqqqqqqqqpmZmZmZmYiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d2ZmZmZmZnd3d3d3d3d3d3d3d3d3d4iIiHd3d4iIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZnd3d2ZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZlVVVVVVVURERFVVVURERERERERERERERDMzM0RERERERDMzM0RERFVVVURERFVVVVVVVWZmZmZmZkRERFVVVVVVVVVVVVVVVURERGZmZmZmZlVVVWZmZnd3d1VVVWZmZoiIiGZmZiIiIiIiIkRERERERFVVVWZmZoiIiJmZmYiIiGZmZlVVVWZmZnd3d2ZmZmZmZmZmZnd3d1VVVURERERERFVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVVVVVURERERERERERERERHd3d5mZmbu7u+7u7szMzIiIiJmZmd3d3bu7u7u7u6qqqqqqqszMzN3d3czMzLu7u6qqqpmZmaqqqszMzMzMzMzMzKqqqpmZmaqqqru7u6qqqoiIiJmZmaqqqru7u7u7u6qqqszMzKqqqpmZmXd3d3d3d4iIiIiIiKqqqpmZmZmZmYiIiHd3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiKqqqpmZmYiIiIiIiJmZmZmZmZmZmYiIiIiIiGZmZnd3d3d3d2ZmZlVVVVVVVWZmZmZmZnd3d3d3d3d3d3d3d2ZmZlVVVVVVVWZmZnd3d4iIiHd3d2ZmZlVVVWZmZmZmZkRERERERFVVVXd3d4iIiHd3d3d3d2ZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZlVVVVVVVXd3d5mZmWZmZkRERGZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZnd3d2ZmZlVVVVVVVVVVVVVVVURERFVVVXd3d2ZmZmZmZlVVVWZmZnd3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZlVVVVVVVXd3d4iIiIiIiIiIiHd3d4iIiHd3d4iIiHd3d2ZmZnd3d3d3d3d3d3d3d4iIiHd3d0RERHd3d6qqqqqqqpmZmXd3d3d3d3d3d4iIiJmZmYiIiHd3d3d3d2ZmZmZmZnd3d2ZmZlVVVWZmZqqqqru7u7u7u6qqqqqqqpmZmZmZmaqqqpmZmaqqqpmZmZmZmaqqqpmZmZmZmYiIiGZmZnd3d5mZmYiIiHd3d3d3d4iIiHd3d3d3d3d3d3d3d4iIiIiIiHd3d4iIiHd3d3d3d3d3d3d3d3d3d4iIiHd3d5mZmbu7u7u7u5mZmYiIiHd3d3d3d2ZmZmZmZmZmZnd3d4iIiIiIiJmZmYiIiGZmZkRERFVVVWZmZmZmZnd3d5mZmaqqqqqqqoiIiHd3d3d3d3d3d3d3d3d3d3d3d6qqqqqqqoiIiIiIiHd3d2ZmZmZmZnd3d2ZmZnd3d3d3d3d3d4iIiIiIiHd3d4iIiHd3d2ZmZmZmZmZmZnd3d3d3d4iIiHd3d3d3d3d3d2ZmZmZmZkRERDMzM1VVVXd3d2ZmZlVVVWZmZkRERFVVVVVVVXd3d1VVVVVVVVVVVWZmZnd3d4iIiHd3d2ZmZnd3d2ZmZkRERFVVVVVVVVVVVURERERERFVVVVVVVURERDMzM0RERERERERERFVVVVVVVWZmZoiIiHd3d3d3d3d3d3d3d1VVVURERDMzM0RERERERFVVVVVVVVVVVVVVVURERERERERERCIiIjMzM0RERFVVVWZmZmZmZnd3d1VVVVVVVWZmZlVVVURERERERERERERERDMzM0RERDMzMzMzM0RERERERERERFVVVVVVVTMzMzMzMzMzM1VVVWZmZmZmZmZmZmZmZkRERERERERERERERERERERERDMzM0RERDMzMyIiIjMzM0RERDMzMzMzM0RERERERDMzM0RERFVVVWZmZlVVVVVVVVVVVVVVVWZmZlVVVURERERERFVVVWZmZlVVVURERERERERERERERERERERERFVVVURERERERDMzM0RERDMzM0RERFVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERDMzM0RERDMzM0RERERERERERERERFVVVTMzM0RERDMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERDMzMxERERERESIiIiIiIjMzMzMzMyIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzM0RERERERFVVVVVVVVVVVURERERERERERERERERERERERFVVVURERERERERERERERDMzMzMzM0RERDMzM0RERERERERERERERFVVVVVVVURERERERERERERERERERFVVVVVVVURERERERERERERERDMzM0RERERERERERDMzM0RERERERERERERERDMzM0RERERERERERFVVVURERDMzMzMzMzMzM0RERERERERERFVVVURERFVVVVVVVWZmZlVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVURERFVVVWZmZnd3d3d3d1VVVTMzMzMzMyIiIlVVVYiIiFVVVURERDMzMyIiIiIiIiIiIlVVVTMzMzMzMyIiIjMzMzMzMzMzM0RERDMzM0RERDMzM0RERERERERERERERERERERERERERERERERERFVVVURERERERERERERERFVVVURERERERERERERERERERFVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERERERFVVVVVVVVVVVURERERERERERFVVVURERERERERERERERDMzM0RERDMzM0RERDMzM0RERDMzMzMzMzMzM0RERDMzMzMzMyIiIiIiIjMzMzMzMzMzM1VVVVVVVURERDMzM0RERFVVVVVVVURERERERDMzM0RERFVVVXd3d3d3d4iIiHd3d0RERERERERERERERGZmZmZmZlVVVURERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERERERFVVVVVVVURERERERFVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVXd3d3d3d3d3d3d3d3d3d4iIiGZmZjMzM0RERGZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZlVVVVVVVVVVVWZmZnd3d2ZmZkRERERERFVVVWZmZmZmZlVVVURERERERERERFVVVURERFVVVURERERERERERFVVVURERFVVVWZmZlVVVVVVVURERERERERERERERERERERERFVVVURERHd3d5mZmXd3d1VVVVVVVWZmZlVVVWZmZoiIiHd3d0RERDMzM3d3d6qqqru7u6qqqqqqqqqqqnd3d3d3d3d3d3d3d3d3d4iIiGZmZmZmZoiIiLu7u8zMzN3d3ZmZmXd3d2ZmZoiIiIiIiGZmZlVVVVVVVWZmZmZmZmZmZoiIiKqqqszMzMzMzJmZmXd3d0RERERERFVVVXd3d2ZmZmZmZmZmZmZmZlVVVVVVVWZmZnd3d5mZmZmZmXd3d1VVVURERERERDMzM0RERHd3d6qqqszMzN3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////u7u7d3d3d3d3d3d3d3d3u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMzd3d3MzMzMzMzMzMy7u7uqqqq7u7vMzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7u7u7uqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqZmZmqqqqZmZmZmZmZmZmZmZmZmZmZmZmIiIiIiIh3d3d3d3dmZmZmZmZmZmZVVVVVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVERERERERERERERERERERVVVVVVVVVVVVmZmZmZmZERERERERVVVVmZmZVVVVERERmZmZmZmZmZmZ3d3d3d3dVVVVmZmZmZmZVVVUzMzMiIiJERERmZmZmZmZ3d3eIiIiqqqqIiIhmZmZmZmZ3d3eZmZmIiIh3d3d3d3dmZmZVVVUzMzNERERVVVVVVVVERERVVVVERERERERVVVVVVVVVVVVERERERERERERVVVVERERVVVV3d3e7u7vd3d2qqqp3d3eqqqrMzMzMzMzMzMyqqqqqqqq7u7u7u7u7u7uqqqqZmZmqqqq7u7vMzMzd3d27u7u7u7uZmZmZmZmqqqqZmZl3d3d3d3e7u7u7u7u7u7u7u7vMzMyqqqqIiIh3d3dmZmZ3d3eIiIiIiIiZmZmIiIiZmZmIiIh3d3eIiIh3d3d3d3eIiIiZmZmZmZmZmZmqqqqqqqqqqqqqqqq7u7uqqqqZmZm7u7uqqqqZmZmIiIh3d3dmZmZVVVVERERVVVVmZmaZmZmZmZl3d3d3d3d3d3dVVVVVVVV3d3eIiIh3d3d3d3d3d3dmZmZVVVVVVVVVVVVERERERERVVVV3d3d3d3d3d3eIiIh3d3d3d3dmZmZ3d3eIiIiIiIh3d3dmZmZmZmZmZmZVVVVmZmZ3d3dmZmZERERmZmaIiIh3d3dmZmZmZmZmZmZVVVVVVVVmZmZmZmZVVVVVVVVEREREREREREQzMzNERERmZmaIiIh3d3d3d3dmZmZmZmZ3d3d3d3d3d3d3d3dmZmZmZmZ3d3dmZmZ3d3d3d3dmZmZ3d3eIiIiIiIiZmZmZmZl3d3eZmZmIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3eIiIiIiIhVVVVmZmaqqqqqqqqqqqqIiIiIiIiIiIiIiIiIiIiZmZl3d3dmZmZ3d3d3d3dmZmZ3d3dmZmZVVVWIiIi7u7vMzMy7u7uZmZmZmZmZmZmZmZmZmZmqqqqqqqqZmZmZmZmIiIh3d3dVVVVVVVVVVVWZmZmZmZl3d3eIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIh3d3eIiIiIiIh3d3eIiIiIiIhmZmZ3d3d3d3eZmZm7u7vMzMy7u7uqqqqIiIh3d3d3d3dmZmZmZmZ3d3eIiIiqqqqZmZl3d3d3d3dmZmZmZmZmZmZmZmZ3d3eIiIiZmZmZmZmIiIh3d3dmZmZ3d3d3d3dmZmaIiIiqqqqZmZmZmZmIiIh3d3dmZmZmZmZVVVVVVVVmZmZmZmZmZmZ3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3d3d3eIiIiIiIiIiIh3d3d3d3d3d3dVVVVERERERERVVVVmZmZVVVVVVVVERERVVVVVVVVVVVVmZmZmZmZERERVVVVmZmZ3d3eIiIh3d3d3d3d3d3d3d3dVVVVERERERERVVVVERERERERVVVVVVVVVVVUzMzMzMzNERERERERVVVVmZmZ3d3eIiIh3d3dmZmZ3d3dmZmZEREREREQzMzNERERERERERERERERERERVVVVVVVVEREREREQzMzMzMzMzMzNmZmZ3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVEREREREQzMzNEREREREQzMzMzMzNERERVVVVVVVVEREREREQzMzMzMzMzMzNVVVVmZmZ3d3dmZmZmZmZVVVVEREREREREREQzMzMzMzMzMzNEREQzMzMzMzMzMzNEREREREREREREREREREQzMzNERERmZmZ3d3dmZmZVVVVVVVVmZmZVVVVmZmZVVVVERERVVVVVVVVERERERERERERERERERERERERERERERERERERERERERERVVVVERERVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVEREREREQzMzMzMzMzMzNEREQzMzNEREREREREREREREREREQzMzMzMzMzMzMzMzNEREREREREREQzMzNEREREREQzMzMREREREREiIiIzMzMzMzMiIiIzMzMzMzMiIiIzMzMiIiIiIiIzMzMiIiIiIiIiIiJERERERERVVVVVVVVVVVVVVVVVVVVEREREREREREREREREREREREREREREREREREQzMzNEREQzMzMzMzNEREREREQzMzNERERERERERERVVVVVVVVERERERERERERVVVVERERERERERERVVVVEREREREREREREREREREREREREREREREQzMzNEREREREREREREREREREREREREREQzMzNERERERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVmZmZ3d3dmZmZmZmZVVVVVVVVVVVVVVVV3d3eIiIh3d3dmZmYzMzMiIiIiIiIzMzOIiIh3d3dmZmYzMzMzMzMiIiIzMzNmZmZEREQzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNEREREREQzMzNERERERERERERERERERERVVVVERERERERERERERERERERERERERERERERERERERERERERERERERERVVVVEREREREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNVVVVVVVVVVVVVVVVEREREREREREREREREREREREREREQzMzNERERERERERERERERERERVVVVEREREREQzMzNEREQzMzMzMzMzMzMiIiIiIiIzMzMzMzNERER3d3dmZmZERERERERERERVVVVVVVVERERERERERERERERVVVV3d3dmZmZmZmZVVVVVVVVEREQzMzNERERmZmZ3d3dmZmZERERVVVUzMzMzMzMzMzMzMzMzMzNEREQzMzNERERERERVVVVERERVVVVVVVVmZmZ3d3dmZmZVVVVVVVVVVVVERERVVVVmZmZ3d3d3d3dmZmZmZmZ3d3d3d3dEREQiIiJERERVVVVmZmZ3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVERERERERmZmaZmZlmZmZERERVVVV3d3d3d3d3d3dVVVVERERERERERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERERERERERVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmYzMzNERER3d3eqqqqqqqqqqqq7u7uqqqpmZmZVVVWIiIiIiIh3d3eIiIh3d3d3d3eZmZm7u7vu7u7u7u7u7u67u7uZmZmZmZmIiIh3d3dVVVVERERERERERERERERmZmZ3d3eIiIiqqqqqqqqIiIhVVVVERERERERVVVVVVVVVVVV3d3dmZmZVVVVVVVVVVVVmZmaIiIiqqqqIiIhmZmZEREQzMzNEREQzMzNERESIiIjMzMzMzMzMzMzu7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u3d3dzMzM3d3d7u7u7u7u3d3d7u7u3d3d7u7u7u7u7u7u3d3d7u7u3d3d7u7u3d3d3d3d3d3d7u7u3d3d7u7u3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMu7u7zMzMu7u7u7u7u7u7u7u7qqqqqqqqmZmZmZmZmZmZiIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3ZmZmd3d3ZmZmVVVVVVVVVVVVREREREREREREREREREREREREREREREREMzMzREREREREREREMzMzREREREREREREREREREREMzMzREREMzMzREREREREREREREREREREREREREREREREREREREREREREREREREREMzMzREREREREREREMzMzREREMzMzREREREREREREREREREREREREREREREREREREVVVVREREREREREREREREVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmd3d3ZmZmZmZmd3d3ZmZmd3d3ZmZmd3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREZmZmVVVVVVVVZmZmd3d3ZmZmd3d3iIiIZmZmVVVVZmZmVVVVMzMzMzMzREREVVVVZmZmd3d3mZmZiIiId3d3d3d3iIiIiIiIiIiIiIiImZmZiIiIVVVVREREREREREREVVVVREREREREVVVVVVVVREREVVVVVVVVREREREREREREREREREREMzMzREREd3d3zMzM3d3dqqqqmZmZqqqqzMzM3d3dzMzMqqqqqqqqqqqqqqqqqqqqqqqqqqqqu7u7zMzM3d3dzMzMqqqqu7u7mZmZiIiImZmZmZmZZmZmiIiIqqqqqqqqu7u7u7u7u7u7qqqqmZmZiIiId3d3iIiIiIiId3d3d3d3iIiImZmZmZmZiIiIiIiIZmZmZmZmmZmZqqqqqqqqqqqqu7u7u7u7qqqqzMzMu7u7qqqqqqqqqqqqqqqqmZmZiIiId3d3ZmZmVVVVVVVVVVVVd3d3mZmZmZmZd3d3ZmZmZmZmVVVVZmZmiIiId3d3d3d3ZmZmd3d3d3d3ZmZmVVVVREREVVVVVVVVVVVVZmZmiIiId3d3iIiIiIiId3d3d3d3d3d3d3d3iIiId3d3ZmZmZmZmZmZmVVVVVVVVVVVVREREREREZmZmiIiId3d3d3d3d3d3ZmZmd3d3ZmZmZmZmZmZmVVVVVVVVREREREREMzMzREREVVVVZmZmiIiId3d3iIiId3d3iIiId3d3iIiId3d3d3d3d3d3ZmZmd3d3d3d3d3d3VVVVVVVVZmZmiIiImZmZmZmZiIiId3d3iIiImZmZiIiIiIiImZmZiIiId3d3ZmZmd3d3d3d3d3d3VVVVZmZmqqqqqqqqqqqqqqqqiIiIiIiIiIiImZmZmZmZiIiId3d3ZmZmVVVVZmZmiIiIZmZmVVVViIiIu7u7u7u7zMzMu7u7u7u7iIiId3d3mZmZqqqqqqqqiIiId3d3ZmZmVVVVVVVVREREVVVVmZmZmZmZmZmZmZmZiIiId3d3iIiIiIiId3d3iIiIiIiId3d3d3d3iIiId3d3iIiId3d3d3d3ZmZmZmZmiIiIqqqqzMzMu7u7qqqqiIiId3d3iIiId3d3d3d3iIiIqqqqmZmZiIiId3d3mZmZiIiId3d3VVVVZmZmZmZmZmZmd3d3iIiIiIiId3d3d3d3d3d3ZmZmd3d3mZmZqqqqmZmZiIiIiIiIiIiId3d3VVVVVVVVZmZmVVVVZmZmd3d3iIiId3d3ZmZmd3d3ZmZmZmZmd3d3ZmZmZmZmiIiImZmZiIiIiIiIiIiIZmZmREREREREREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmd3d3d3d3iIiIiIiId3d3d3d3ZmZmVVVVVVVVVVVVREREVVVVREREREREVVVVREREREREMzMzIiIiMzMzREREd3d3iIiIiIiId3d3ZmZmZmZmZmZmVVVVMzMzREREREREREREREREVVVVREREVVVVVVVVREREREREMzMzREREREREZmZmd3d3ZmZmd3d3ZmZmVVVVVVVVREREVVVVREREREREREREREREREREREREMzMzREREVVVVREREREREMzMzMzMzIiIiMzMzVVVVZmZmZmZmZmZmVVVVVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREIiIiMzMzZmZmd3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREMzMzMzMzREREREREREREVVVVREREMzMzMzMzVVVVZmZmVVVVZmZmZmZmZmZmZmZmVVVVVVVVREREVVVVREREREREREREMzMzREREMzMzMzMzREREREREREREREREREREMzMzMzMzMzMzREREREREREREVVVVMzMzMzMzREREMzMzERERIiIiIiIiMzMzMzMzMzMzIiIiMzMzIiIiIiIiMzMzIiIiIiIiIiIiIiIiMzMzVVVVREREREREVVVVVVVVVVVVZmZmVVVVREREVVVVREREVVVVREREREREREREMzMzREREREREREREMzMzMzMzREREREREREREVVVVREREREREVVVVREREREREVVVVREREREREVVVVREREREREREREREREREREREREVVVVREREREREMzMzMzMzMzMzMzMzREREREREREREREREREREMzMzMzMzMzMzREREVVVVZmZmREREVVVVVVVVZmZmVVVVVVVVVVVVZmZmZmZmVVVVVVVVREREZmZmd3d3iIiIZmZmVVVVVVVVVVVVVVVVd3d3iIiImZmZiIiIZmZmMzMzMzMzIiIiMzMzmZmZiIiIVVVVREREIiIiIiIiMzMzVVVVVVVVMzMzIiIiIiIiIiIiMzMzMzMzREREREREREREREREREREMzMzREREREREREREVVVVVVVVREREREREREREREREREREREREREREREREREREREREVVVVREREVVVVVVVVVVVVREREREREREREMzMzREREMzMzMzMzMzMzMzMzREREMzMzVVVVd3d3ZmZmREREVVVVREREREREREREREREREREREREMzMzREREMzMzREREREREREREVVVVZmZmVVVVMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzREREd3d3ZmZmREREREREREREVVVVVVVVZmZmVVVVREREREREVVVViIiId3d3VVVVVVVVVVVVREREREREVVVVZmZmd3d3iIiIVVVVREREMzMzMzMzMzMzREREMzMzMzMzMzMzREREVVVVVVVVREREVVVVd3d3d3d3d3d3iIiIZmZmREREREREREREVVVVVVVVd3d3d3d3ZmZmZmZmd3d3iIiIVVVVMzMzMzMzREREZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREVVVVmZmZiIiIREREREREZmZmZmZmVVVVREREREREMzMzREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREMzMzREREREREREREREREREREVVVVVVVVREREREREVVVVVVVVVVVVVVVVVVVVZmZmVVVVMzMzVVVVd3d3mZmZqqqqzMzMu7u7iIiIVVVVd3d3iIiIiIiIiIiIiIiId3d3iIiIqqqqu7u73d3d7u7u3d3d3d3du7u7qqqqmZmZmZmZmZmZd3d3VVVVREREVVVVVVVVd3d3ZmZmZmZmd3d3ZmZmREREVVVVREREREREVVVVREREVVVVZmZmZmZmVVVVVVVVZmZmZmZmiIiImZmZiIiIVVVVREREREREMzMzREREd3d3qqqqzMzMu7u7zMzM3d3d////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////+7u7t3d3d3d3d3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3e7u7t3d3e7u7t3d3d3d3e7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzLu7u7u7u7u7u6qqqqqqqqqqqpmZmZmZmZmZmZmZmXd3d4iIiHd3d3d3d2ZmZmZmZmZmZkRERFVVVVVVVVVVVURERERERERERERERFVVVURERERERERERERERERERERERERERERERDMzM0RERERERERERDMzMzMzMzMzM0RERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERDMzMzMzM0RERDMzM0RERERERERERFVVVWZmZlVVVWZmZmZmZmZmZmZmZnd3d2ZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZlVVVWZmZlVVVVVVVWZmZnd3d2ZmZmZmZnd3d1VVVVVVVWZmZlVVVTMzMzMzM0RERFVVVWZmZnd3d4iIiIiIiIiIiIiIiHd3d3d3d3d3d4iIiKqqqoiIiFVVVURERERERFVVVVVVVURERFVVVURERERERERERFVVVVVVVURERERERERERERERERERCIiIkRERHd3d6qqqt3d3aqqqru7u7u7u7u7u7u7u8zMzKqqqpmZmbu7u6qqqqqqqqqqqru7u93d3d3d3czMzLu7u6qqqpmZmZmZmZmZmZmZmZmZmXd3d3d3d5mZmaqqqru7u7u7u7u7u6qqqqqqqqqqqpmZmZmZmZmZmYiIiIiIiHd3d3d3d4iIiJmZmXd3d1VVVWZmZpmZmbu7u7u7u6qqqqqqqqqqqru7u8zMzLu7u6qqqqqqqqqqqqqqqpmZmYiIiHd3d3d3d4iIiGZmZlVVVWZmZpmZmaqqqoiIiGZmZnd3d2ZmZoiIiIiIiHd3d3d3d4iIiHd3d3d3d4iIiHd3d0RERERERERERFVVVXd3d5mZmXd3d3d3d4iIiJmZmXd3d3d3d3d3d4iIiHd3d3d3d3d3d2ZmZmZmZmZmZkRERERERERERHd3d5mZmYiIiIiIiHd3d4iIiHd3d3d3d2ZmZmZmZmZmZlVVVURERERERERERERERFVVVWZmZnd3d3d3d3d3d4iIiIiIiIiIiIiIiHd3d4iIiIiIiHd3d2ZmZnd3d2ZmZlVVVURERFVVVZmZmZmZmYiIiJmZmYiIiIiIiIiIiHd3d4iIiJmZmZmZmXd3d2ZmZmZmZnd3d2ZmZlVVVWZmZpmZmaqqqqqqqqqqqoiIiIiIiIiIiJmZmZmZmZmZmXd3d2ZmZmZmZnd3d3d3d3d3d2ZmZoiIiMzMzLu7u8zMzMzMzLu7u6qqqqqqqqqqqpmZmYiIiGZmZmZmZlVVVVVVVURERERERFVVVXd3d6qqqpmZmZmZmXd3d3d3d4iIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d5mZmYiIiIiIiHd3d1VVVVVVVWZmZnd3d6qqqru7u6qqqoiIiIiIiIiIiJmZmYiIiHd3d5mZmYiIiHd3d5mZmZmZmXd3d2ZmZlVVVVVVVWZmZlVVVXd3d5mZmaqqqoiIiHd3d2ZmZmZmZoiIiKqqqpmZmYiIiJmZmZmZmYiIiHd3d1VVVVVVVVVVVVVVVWZmZmZmZoiIiHd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZoiIiJmZmYiIiIiIiGZmZmZmZlVVVURERERERGZmZmZmZkRERFVVVVVVVVVVVVVVVURERFVVVVVVVVVVVWZmZoiIiIiIiIiIiHd3d4iIiIiIiGZmZlVVVVVVVURERERERERERERERERERFVVVURERERERDMzMzMzMyIiIlVVVYiIiIiIiHd3d3d3d1VVVWZmZlVVVVVVVVVVVURERERERFVVVURERERERERERFVVVVVVVURERERERERERERERFVVVWZmZmZmZmZmZnd3d2ZmZlVVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERERERFVVVURERERERDMzMyIiIjMzM0RERFVVVWZmZmZmZmZmZlVVVURERERERERERERERERERDMzMzMzMzMzMzMzMzMzMyIiIjMzM0RERDMzMzMzMyIiIjMzMzMzM1VVVWZmZmZmZmZmZmZmZlVVVURERFVVVVVVVURERERERERERERERDMzMzMzM0RERDMzM0RERFVVVURERERERDMzM1VVVWZmZlVVVWZmZnd3d2ZmZmZmZlVVVWZmZlVVVVVVVVVVVURERDMzM0RERDMzM0RERDMzMzMzM0RERERERERERERERERERDMzMzMzM0RERERERERERERERERERERERERERDMzMxERESIiIiIiIkRERERERDMzMzMzMyIiIjMzMyIiIiIiIjMzMyIiIiIiIjMzMzMzM1VVVVVVVVVVVURERGZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERERERDMzM0RERDMzMzMzM0RERFVVVVVVVVVVVURERERERERERFVVVURERERERFVVVURERERERERERERERFVVVVVVVWZmZkRERERERERERERERDMzM0RERDMzM0RERERERERERDMzMzMzMzMzM0RERHd3d1VVVURERFVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVURERFVVVURERHd3d5mZmZmZmVVVVVVVVWZmZlVVVVVVVWZmZnd3d3d3d3d3d1VVVTMzMzMzMyIiIjMzM4iIiJmZmWZmZkRERDMzMzMzMyIiIlVVVWZmZjMzMxERESIiIjMzM0RERDMzMzMzM0RERERERDMzM0RERERERDMzM0RERERERERERERERERERERERERERERERERERERERERERERERERERERERFVVVVVVVURERGZmZmZmZkRERERERERERDMzMzMzMzMzM0RERERERERERERERERERFVVVXd3d2ZmZkRERERERERERERERERERERERERERDMzM0RERDMzMzMzM0RERFVVVVVVVWZmZmZmZkRERDMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERDMzM0RERFVVVWZmZlVVVURERERERFVVVVVVVVVVVWZmZlVVVVVVVWZmZnd3d3d3d1VVVURERFVVVURERERERFVVVVVVVXd3d4iIiFVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVURERGZmZnd3d2ZmZnd3d3d3d1VVVVVVVURERERERGZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3dzMzMzMzM0RERFVVVWZmZnd3d2ZmZlVVVVVVVVVVVVVVVVVVVURERFVVVURERERERFVVVYiIiKqqqpmZmWZmZkRERERERFVVVURERERERGZmZmZmZkRERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERERERFVVVVVVVURERFVVVURERERERERERERERERERFVVVURERFVVVVVVVVVVVWZmZlVVVTMzM1VVVYiIiLu7u7u7u6qqqoiIiGZmZmZmZnd3d4iIiHd3d2ZmZnd3d4iIiJmZmczMzLu7u7u7u8zMzMzMzN3d3czMzKqqqqqqqszMzMzMzKqqqnd3d1VVVURERFVVVXd3d2ZmZlVVVVVVVURERERERERERERERDMzM0RERDMzM0RERFVVVVVVVWZmZlVVVWZmZmZmZnd3d3d3d4iIiIiIiFVVVURERERERDMzM1VVVZmZmbu7u8zMzKqqqru7u+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////d3d3u7u7u7u7u7u7////u7u7////u7u7u7u7u7u7u7u7d3d3d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3MzMzd3d3d3d3d3d3d3d3u7u7d3d3u7u7d3d3u7u7d3d3u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7u7u7d3d3d3d3u7u7d3d3u7u7d3d3d3d3d3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMy7u7u7u7uqqqqqqqqqqqqqqqqZmZmqqqqIiIiIiIiIiIiIiIh3d3d3d3eIiIh3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVEREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNEREQzMzMzMzNEREQzMzMzMzMzMzNEREREREQzMzMzMzMzMzNEREREREREREQzMzNEREREREREREQzMzNERERERERERERERERERERVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZ3d3d3d3dmZmZ3d3d3d3d3d3d3d3dmZmZ3d3dmZmZVVVVVVVVVVVVmZmZVVVVERERVVVVVVVVmZmZ3d3dERERVVVVmZmZVVVV3d3eIiIh3d3eZmZmZmZl3d3dVVVVVVVVmZmZmZmZ3d3d3d3dVVVVERERVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVEREREREQzMzMzMzNEREREREQzMzNERERmZmaIiIi7u7u7u7vMzMzMzMy7u7u7u7u7u7uqqqqZmZmqqqqqqqqqqqrMzMzMzMzMzMzd3d3MzMzMzMyqqqqqqqqqqqqqqqq7u7uqqqqIiIh3d3d3d3eZmZmqqqq7u7u7u7u7u7u7u7u7u7u7u7uZmZmZmZmZmZmIiIhmZmaIiIiIiIiIiIh3d3dmZmZmZmaIiIi7u7u7u7uqqqq7u7u7u7u7u7u7u7vMzMy7u7uqqqqqqqqZmZmZmZmIiIh3d3eIiIi7u7t3d3dVVVV3d3eqqqqqqqqIiIh3d3dmZmaIiIiZmZmIiIiIiIiIiIiZmZmZmZmIiIh3d3dmZmZERERERERVVVVmZmaIiIiIiIiIiIh3d3eIiIiZmZmIiIh3d3d3d3eIiIiIiIiIiIiIiIh3d3d3d3dmZmZmZmZmZmZmZmZ3d3eqqqqZmZl3d3d3d3d3d3eIiIh3d3dmZmZmZmZ3d3dmZmZmZmZVVVVERERERERmZmZ3d3eIiIiIiIh3d3eIiIiZmZmZmZmZmZmIiIiIiIiIiIh3d3d3d3dmZmZ3d3d3d3dVVVVVVVWIiIiZmZmZmZmqqqqIiIiIiIiIiIiIiIiIiIh3d3eIiIiIiIh3d3d3d3dmZmZmZmZVVVVmZmaqqqqqqqqqqqqZmZmIiIiqqqqZmZmIiIiZmZmIiIh3d3dmZmZ3d3eZmZmIiIhmZmZmZmaZmZnMzMzMzMy7u7u7u7vMzMzMzMy7u7uqqqqIiIhmZmZVVVVVVVVVVVVERERVVVVVVVVmZmaIiIiZmZmZmZmZmZmZmZmIiIiIiIiIiIh3d3d3d3eIiIh3d3d3d3eIiIiZmZmZmZmIiIh3d3dmZmZmZmZERERVVVWIiIi7u7uqqqqZmZmIiIiZmZmZmZmIiIh3d3eIiIiZmZmZmZmqqqp3d3dmZmZERERERERVVVVmZmZ3d3d3d3eZmZmZmZl3d3dmZmZVVVVmZmaIiIiZmZmqqqqqqqqqqqqZmZl3d3dVVVVVVVVVVVVERERVVVVmZmZmZmaIiIhmZmZmZmZmZmZmZmZ3d3dmZmZmZmZ3d3eIiIiZmZmIiIh3d3dVVVVVVVVmZmZVVVVVVVVmZmZVVVVVVVVVVVVERERERERVVVVEREQzMzNERERERERmZmaIiIiZmZl3d3dmZmZ3d3dmZmZVVVVVVVVVVVVERERERERERERERERERERVVVVVVVVEREQzMzMiIiIzMzNVVVWIiIiZmZl3d3dVVVVmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVmZmZ3d3dmZmZ3d3d3d3dmZmZmZmZERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERVVVVEREQzMzNEREQzMzNERERVVVVmZmZmZmZmZmZVVVVVVVVVVVVEREREREREREREREQzMzMzMzMiIiIzMzMzMzMzMzMzMzNEREQzMzMzMzMiIiIzMzMzMzNVVVVmZmZmZmZmZmZVVVVERERVVVVEREREREREREREREREREREREREREQzMzNEREQzMzNEREQzMzNEREREREQzMzNERERVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVmZmZVVVVEREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzNEREREREQzMzMzMzMzMzMzMzNVVVVVVVUzMzMiIiIiIiIREREzMzMzMzMzMzMzMzMiIiIiIiIiIiIzMzMzMzMzMzMzMzMiIiJERERERERVVVVERERVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVEREREREREREQzMzNEREREREREREQzMzMzMzNERERVVVVERERERERERERVVVVERERERERERERERERERERERERERERVVVVVVVVmZmZmZmZVVVVVVVVEREREREREREREREQzMzNEREREREREREREREQzMzMzMzNVVVV3d3dVVVVERERERERVVVVVVVVVVVVVVVVERERERERERERERERERERmZmaZmZmqqqpmZmZERERmZmZmZmZmZmZmZmZ3d3dmZmZmZmZVVVVEREQzMzMzMzMzMzMzMzN3d3eqqqp3d3dEREREREREREREREREREREREQiIiIREREzMzMzMzNEREQzMzNEREREREQzMzNEREREREQzMzMzMzNERERERERERERERERERERERERERERERERERERERERERERERERERERVVVVERERERERERERVVVVVVVUzMzMzMzMzMzMzMzNERERERERERERVVVVVVVVERERVVVVVVVVmZmZEREQzMzMzMzNEREREREREREREREREREQzMzMzMzNEREQzMzNERERERERmZmZVVVVVVVUzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVVVVVERERVVVVVVVVmZmZVVVVVVVVmZmZVVVVmZmZmZmZVVVUzMzNERERERERERERVVVVERERVVVVVVVV3d3dmZmZEREREREREREQzMzMzMzMzMzMzMzMzMzNERERERERERERERERmZmZmZmZmZmZmZmZ3d3dVVVVVVVVVVVVmZmZ3d3dmZmZmZmZ3d3dmZmZVVVVmZmZ3d3d3d3dVVVUzMzMzMzNERERmZmZmZmZ3d3dVVVVERERVVVVERERVVVVERERVVVVERERERERERERVVVV3d3fMzMy7u7tmZmZEREQzMzMzMzNmZmaIiIh3d3dVVVVERERmZmZVVVVERERVVVVERERERERERERERERERERERERERERERERVVVVERERmZmZVVVVERERERERVVVVVVVVVVVVVVVVVVVVERERVVVVmZmZVVVUzMzNERER3d3eZmZm7u7uZmZl3d3dmZmZmZmaIiIiIiIhmZmZmZmZmZmZ3d3eIiIiqqqqqqqqqqqqIiIiIiIjMzMzu7u7u7u7u7u7d3d3MzMyqqqqZmZl3d3dVVVVERERERERmZmZ3d3dmZmZVVVVEREREREQzMzNEREREREQzMzMzMzMzMzMzMzNERERVVVVVVVVmZmZ3d3d3d3dmZmZ3d3d3d3dmZmZVVVUzMzNERERERERVVVWqqqrMzMy7u7uqqqrMzMzu7u7u7u7////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u7u7u3d3d3d3d7u7u3d3d7u7u3d3d3d3d3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d7u7u7u7u3d3d7u7u7u7u7u7u7u7u3d3d7u7u3d3d7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMu7u7zMzMu7u7u7u7u7u7u7u7u7u7u7u7qqqqu7u7u7u7u7u7qqqqqqqqqqqqqqqqmZmZmZmZqqqqmZmZmZmZiIiImZmZiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3d3d3ZmZmVVVVVVVVREREVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzREREREREREREMzMzREREREREVVVVREREVVVVVVVVVVVVZmZmZmZmREREREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVREREREREREREREREVVVVREREREREREREVVVVVVVVVVVVVVVVZmZmd3d3d3d3ZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmd3d3VVVVZmZmZmZmZmZmiIiIiIiId3d3iIiImZmZZmZmREREREREVVVVVVVVVVVVZmZmREREREREREREREREREREVVVVZmZmVVVVVVVVVVVVREREMzMzREREREREMzMzVVVVVVVVMzMzREREREREZmZmqqqqu7u7u7u7u7u7zMzMzMzMzMzMu7u7iIiIqqqqqqqqu7u73d3dzMzMu7u7u7u7u7u7u7u7zMzMu7u7u7u7u7u7qqqqqqqqiIiId3d3ZmZmqqqqu7u7qqqqqqqqqqqqu7u7u7u7qqqqiIiIiIiImZmZiIiIiIiIiIiImZmZiIiIiIiId3d3ZmZmZmZmiIiIu7u7u7u7u7u7zMzMu7u7u7u7zMzMzMzMu7u7mZmZqqqqmZmZiIiId3d3iIiImZmZiIiIZmZmiIiIqqqqqqqqiIiIiIiIiIiIiIiIqqqqqqqqmZmZiIiImZmZqqqqmZmZd3d3ZmZmVVVVREREVVVViIiImZmZqqqqmZmZiIiImZmZiIiIiIiImZmZmZmZiIiIiIiImZmZmZmZd3d3d3d3ZmZmVVVVZmZmd3d3mZmZiIiIiIiIiIiId3d3iIiIiIiIiIiId3d3ZmZmZmZmZmZmd3d3VVVVREREREREd3d3d3d3iIiId3d3mZmZqqqqmZmZqqqqmZmZmZmZiIiIiIiId3d3d3d3ZmZmZmZmiIiIZmZmREREd3d3qqqqmZmZqqqqmZmZiIiIiIiIiIiIiIiImZmZiIiId3d3d3d3d3d3ZmZmZmZmZmZmZmZmmZmZu7u7qqqqqqqqmZmZqqqqqqqqmZmZmZmZiIiId3d3ZmZmiIiImZmZmZmZd3d3VVVViIiIu7u73d3du7u7zMzMzMzMzMzMqqqqd3d3ZmZmZmZmVVVVREREVVVVVVVVVVVVVVVVZmZmd3d3iIiIqqqqqqqqmZmZiIiIiIiId3d3d3d3d3d3iIiId3d3d3d3qqqqmZmZiIiIiIiIZmZmZmZmZmZmREREREREVVVVqqqqu7u7mZmZmZmZmZmZiIiIZmZmZmZmqqqqu7u7qqqqiIiIZmZmVVVVVVVVVVVVVVVVZmZmd3d3d3d3d3d3mZmZd3d3d3d3ZmZmZmZmd3d3mZmZqqqqqqqqqqqqiIiId3d3VVVVREREREREVVVVREREVVVVZmZmiIiIZmZmZmZmZmZmZmZmZmZmZmZmZmZmiIiIiIiImZmZiIiIiIiIZmZmVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREREREREREMzMzREREREREZmZmmZmZiIiId3d3ZmZmZmZmZmZmZmZmVVVVREREMzMzREREREREREREREREVVVVVVVVVVVVMzMzMzMzIiIiZmZmiIiIiIiIiIiId3d3ZmZmZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVREREVVVVREREVVVVVVVVVVVVd3d3ZmZmZmZmZmZmd3d3VVVVVVVVVVVVVVVVVVVVREREREREVVVVVVVVVVVVREREREREREREREREREREREREREREMzMzREREVVVVVVVVZmZmZmZmVVVVVVVVREREREREREREMzMzREREREREREREMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVREREREREREREMzMzREREREREREREREREMzMzREREREREREREREREREREVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVREREMzMzREREREREMzMzMzMzMzMzREREREREREREIiIiMzMzREREREREMzMzMzMzMzMzREREZmZmREREIiIiIiIiIiIiERERIiIiIiIiIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzIiIiREREVVVVVVVVVVVVREREZmZmZmZmZmZmZmZmREREREREREREREREREREREREVVVVREREREREREREREREREREREREREREMzMzMzMzREREREREREREREREVVVVREREVVVVREREVVVVREREREREREREREREVVVVZmZmZmZmZmZmVVVVVVVVREREREREREREREREMzMzREREREREREREREREREREMzMzREREZmZmVVVVREREVVVVVVVVREREVVVVREREVVVVVVVVVVVVVVVVREREd3d3qqqqiIiIZmZmREREVVVVd3d3ZmZmd3d3d3d3ZmZmZmZmVVVVVVVVREREMzMzREREMzMzd3d3qqqqmZmZZmZmVVVVREREREREREREIiIiERERIiIiIiIiREREMzMzMzMzMzMzMzMzREREMzMzMzMzREREREREREREMzMzMzMzREREMzMzREREREREREREREREREREMzMzREREREREVVVVREREREREREREREREVVVVREREMzMzMzMzMzMzVVVVREREVVVVZmZmVVVVREREREREVVVVVVVVREREREREREREMzMzREREREREREREMzMzREREREREMzMzREREREREZmZmZmZmVVVVREREMzMzMzMzIiIiMzMzREREREREMzMzMzMzREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVREREVVVVVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVVVVVVVVVVVVVZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmVVVVZmZmZmZmREREMzMzMzMzREREZmZmZmZmVVVVVVVVREREREREVVVVVVVVVVVVVVVVREREREREMzMzREREmZmZzMzMqqqqVVVVREREMzMzREREZmZmREREMzMzZmZmd3d3ZmZmVVVVREREREREREREREREREREREREREREREREREREREREVVVVREREVVVVVVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVViIiIqqqqqqqqd3d3ZmZmZmZmiIiIqqqqmZmZZmZmZmZmZmZmZmZmd3d3d3d3iIiIqqqqqqqqmZmZ3d3d7u7u7u7u3d3du7u7mZmZd3d3d3d3d3d3VVVVVVVVREREVVVVVVVVZmZmVVVVVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREVVVVVVVVZmZmd3d3d3d3ZmZmVVVVZmZmVVVVREREREREREREVVVVd3d3u7u7zMzMqqqqzMzM7u7u7u7u////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////+7u7v///////////////////////////////+7u7t3d3e7u7u7u7u7u7u7u7u7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7u7u7t3d3e7u7u7u7t3d3e7u7u7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3e7u7t3d3d3d3d3d3czMzN3d3d3d3czMzMzMzMzMzN3d3czMzMzMzMzMzMzMzMzMzMzMzLu7u7u7u8zMzLu7u7u7u6qqqru7u7u7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqru7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqpmZmZmZmaqqqpmZmZmZmYiIiHd3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVURERERERFVVVURERERERDMzM0RERERERERERERERERERFVVVURERERERERERERERDMzM0RERERERERERFVVVVVVVURERFVVVVVVVVVVVWZmZlVVVWZmZnd3d2ZmZmZmZlVVVVVVVVVVVWZmZnd3d2ZmZmZmZnd3d3d3d2ZmZlVVVVVVVURERFVVVVVVVVVVVVVVVURERFVVVWZmZlVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d2ZmZnd3d4iIiHd3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiHd3d2ZmZlVVVVVVVURERERERFVVVURERFVVVURERERERDMzM0RERGZmZnd3d2ZmZlVVVVVVVURERERERERERERERERERERERERERDMzM0RERERERGZmZqqqqru7u7u7u7u7u8zMzN3d3d3d3aqqqnd3d6qqqru7u8zMzN3d3d3d3bu7u7u7u6qqqqqqqru7u7u7u7u7u7u7u7u7u6qqqpmZmXd3d4iIiLu7u6qqqqqqqqqqqszMzMzMzMzMzJmZmZmZmZmZmYiIiIiIiIiIiIiIiHd3d3d3d4iIiHd3d1VVVXd3d4iIiMzMzMzMzLu7u7u7u8zMzMzMzMzMzMzMzLu7u6qqqqqqqqqqqoiIiHd3d3d3d4iIiIiIiHd3d5mZmaqqqqqqqru7u6qqqqqqqpmZmaqqqru7u5mZmYiIiJmZmZmZmYiIiHd3d2ZmZlVVVVVVVWZmZoiIiKqqqru7u6qqqpmZmZmZmZmZmZmZmZmZmaqqqqqqqpmZmYiIiIiIiIiIiIiIiHd3d2ZmZlVVVYiIiJmZmYiIiIiIiIiIiIiIiJmZmYiIiHd3d3d3d2ZmZlVVVXd3d3d3d1VVVVVVVURERFVVVXd3d4iIiIiIiIiIiJmZmaqqqpmZmaqqqpmZmZmZmYiIiHd3d3d3d3d3d2ZmZnd3d2ZmZlVVVXd3d6qqqru7u6qqqqqqqpmZmZmZmYiIiJmZmYiIiIiIiIiIiGZmZnd3d3d3d2ZmZmZmZmZmZqqqqru7u7u7u6qqqpmZmaqqqqqqqoiIiHd3d4iIiJmZmYiIiIiIiIiIiHd3d2ZmZmZmZnd3d6qqqt3d3czMzMzMzLu7u7u7u2ZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVXd3d4iIiKqqqqqqqqqqqpmZmYiIiIiIiHd3d4iIiHd3d3d3d4iIiKqqqoiIiHd3d3d3d3d3d2ZmZlVVVTMzMzMzMzMzM4iIiLu7u6qqqpmZmZmZmXd3d1VVVXd3d6qqqszMzKqqqnd3d2ZmZlVVVVVVVWZmZlVVVWZmZoiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d5mZmbu7u6qqqpmZmXd3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZoiIiHd3d1VVVVVVVVVVVVVVVWZmZlVVVYiIiJmZmZmZmYiIiHd3d3d3d2ZmZlVVVURERFVVVVVVVVVVVVVVVWZmZlVVVVVVVURERFVVVURERERERGZmZnd3d4iIiIiIiIiIiGZmZnd3d2ZmZmZmZkRERERERDMzMzMzMzMzMzMzM0RERERERFVVVURERERERDMzMzMzM3d3d4iIiIiIiHd3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZkRERERERFVVVURERERERFVVVVVVVVVVVVVVVVVVVXd3d2ZmZmZmZmZmZlVVVWZmZlVVVVVVVURERERERFVVVURERFVVVVVVVVVVVURERERERERERERERERERERERERERDMzM1VVVVVVVVVVVVVVVVVVVVVVVURERERERERERDMzMzMzMzMzM0RERERERERERDMzMzMzMzMzMzMzM0RERDMzMyIiIiIiIjMzM1VVVWZmZnd3d1VVVVVVVVVVVVVVVURERERERERERERERFVVVVVVVVVVVURERFVVVURERERERERERERERERERERERERERERERFVVVVVVVWZmZmZmZmZmZmZmZkRERERERERERERERFVVVVVVVVVVVURERERERDMzMzMzM0RERDMzM0RERERERERERCIiIjMzM0RERDMzMzMzMzMzMyIiIjMzM3d3d0RERDMzMyIiIhERESIiIiIiIhERESIiIjMzMyIiIiIiIhERESIiIiIiIiIiIhERESIiIiIiIlVVVXd3d1VVVVVVVVVVVVVVVWZmZlVVVURERERERERERERERFVVVVVVVURERFVVVURERERERERERERERERERERERERERDMzM0RERERERERERDMzM0RERERERFVVVURERFVVVVVVVURERFVVVURERERERFVVVXd3d3d3d2ZmZlVVVVVVVURERERERERERDMzM0RERERERERERFVVVURERERERERERERERERERERERFVVVURERERERFVVVURERFVVVWZmZlVVVVVVVVVVVXd3d6qqqpmZmWZmZlVVVURERFVVVXd3d4iIiIiIiIiIiGZmZlVVVWZmZlVVVURERERERERERDMzM3d3d6qqqpmZmWZmZkRERDMzM1VVVVVVVSIiIhERESIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERDMzM0RERERERERERERERERERERERERERERERERERDMzM0RERERERFVVVURERERERERERDMzM1VVVURERERERDMzM0RERFVVVURERERERFVVVVVVVURERFVVVVVVVURERERERERERDMzM0RERDMzM0RERERERDMzM0RERDMzM0RERERERGZmZnd3d2ZmZlVVVURERDMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzM0RERERERERERERERFVVVVVVVVVVVWZmZmZmZlVVVVVVVURERFVVVVVVVVVVVURERFVVVWZmZlVVVURERERERGZmZmZmZkRERFVVVXd3d3d3d0RERDMzMzMzM0RERERERERERERERFVVVURERFVVVVVVVVVVVVVVVURERFVVVVVVVWZmZnd3d2ZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZlVVVURERCIiIjMzM1VVVWZmZlVVVURERERERFVVVURERFVVVVVVVVVVVURERERERERERDMzM1VVVaqqqszMzGZmZlVVVVVVVTMzMzMzMzMzM2ZmZoiIiIiIiJmZmXd3d1VVVURERERERERERERERERERDMzM0RERERERERERFVVVURERERERERERERERFVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVTMzM0RERHd3d5mZmZmZmXd3d2ZmZmZmZnd3d3d3d6qqqpmZmXd3d2ZmZmZmZlVVVVVVVWZmZoiIiMzMzLu7u6qqqszMzO7u7szMzKqqqoiIiGZmZmZmZmZmZlVVVVVVVVVVVURERFVVVVVVVVVVVWZmZmZmZlVVVURERDMzM0RERDMzMzMzMzMzM0RERDMzM0RERERERERERGZmZnd3d3d3d2ZmZlVVVVVVVURERERERDMzMzMzM0RERFVVVYiIiLu7u8zMzLu7u8zMzN3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7d3d3d3d3u7u7u7u7u7u7u7u7d3d3d3d3d3d3u7u7u7u7d3d3u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3d3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzd3d3MzMzMzMzMzMzMzMy7u7vMzMy7u7vMzMy7u7u7u7u7u7u7u7uqqqqqqqqqqqqZmZmZmZmqqqqZmZmqqqqqqqq7u7uqqqqqqqqqqqq7u7uqqqq7u7u7u7uqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqZmZmqqqqZmZmZmZmZmZmZmZmIiIiIiIiIiIh3d3d3d3d3d3dmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVERERERERERERVVVVERERERERVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVERERVVVVVVVVVVVVmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3dVVVVVVVVVVVVmZmZVVVVVVVV3d3d3d3d3d3dmZmZmZmZmZmZ3d3dmZmZ3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3dmZmZmZmZ3d3d3d3dmZmZ3d3eIiIiIiIiIiIiIiIiIiIhmZmZVVVVVVVVVVVVVVVVmZmZmZmZVVVVERERERERERERVVVVmZmZ3d3dmZmZmZmZERERERERVVVVVVVVVVVVEREQzMzMzMzNERERERERERESIiIiqqqrMzMy7u7uqqqqqqqq7u7uqqqqIiIh3d3eZmZmqqqrMzMzd3d3d3d3d3d27u7u7u7uqqqq7u7vMzMy7u7u7u7u7u7uZmZmIiIiZmZmqqqrMzMyqqqqqqqqqqqq7u7vMzMzMzMy7u7uqqqqZmZmZmZmZmZmIiIh3d3dmZmaIiIiZmZlmZmZmZmZ3d3eZmZnMzMzMzMy7u7u7u7vMzMzMzMzd3d3MzMy7u7u7u7uqqqqZmZl3d3d3d3eIiIh3d3d3d3eIiIiqqqrMzMy7u7u7u7u7u7u7u7vMzMy7u7vMzMyqqqqIiIiIiIiIiIiIiIh3d3d3d3d3d3dVVVV3d3eZmZmqqqq7u7u7u7uqqqqqqqqqqqqqqqqIiIiIiIiZmZmqqqqZmZmZmZmZmZmIiIiIiIh3d3dVVVV3d3eZmZmZmZmZmZmZmZmqqqqZmZmIiIiIiIh3d3dmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVV3d3eIiIiZmZmIiIiIiIiZmZmqqqqZmZmZmZmZmZmIiIiIiIh3d3d3d3dmZmZ3d3dmZmZVVVWIiIiqqqq7u7uqqqq7u7uqqqqqqqqqqqqZmZmIiIiIiIh3d3eIiIh3d3d3d3dmZmZVVVVVVVWIiIi7u7u7u7u7u7uqqqqqqqqZmZl3d3eIiIiIiIiZmZmZmZmIiIh3d3dmZmZ3d3d3d3d3d3eZmZm7u7vMzMzMzMy7u7uIiIhVVVVERERERERVVVVmZmZVVVVmZmZVVVVVVVVERERVVVVmZmaZmZmqqqqqqqqqqqqZmZl3d3d3d3d3d3d3d3d3d3d3d3eqqqqZmZl3d3d3d3dmZmZVVVVEREREREQzMzMzMzNERERVVVWIiIiqqqq7u7uqqqqIiIh3d3eZmZm7u7u7u7uZmZlmZmZVVVVVVVVERERVVVVVVVV3d3eIiIiZmZl3d3dVVVVVVVVmZmaIiIiIiIh3d3eIiIiqqqqZmZmZmZl3d3dVVVVmZmZmZmZVVVVVVVVVVVVVVVVmZmZ3d3dmZmZVVVVmZmZVVVVmZmZVVVVVVVWIiIiZmZmIiIiIiIh3d3dmZmZVVVVVVVVEREREREQzMzNERERVVVVmZmZmZmZVVVVVVVVVVVVERERERERmZmaIiIiqqqqqqqqIiIh3d3d3d3dVVVVVVVVEREREREREREQzMzNEREQzMzNERERVVVVEREREREQzMzMzMzMzMzN3d3eIiIiIiIh3d3dmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZVVVVERERVVVVERERERERERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3dmZmZERERVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVEREREREQzMzNVVVVEREQzMzNERERERERERERmZmZVVVVVVVVERERVVVVEREREREREREREREREREREREREREQzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzNVVVVVVVV3d3d3d3dmZmZmZmZVVVVVVVVERERERERERERERERVVVVVVVVVVVVVVVVEREQzMzMzMzNERERERERERERVVVVVVVVERERVVVVVVVVmZmZ3d3dmZmZVVVVVVVVEREREREREREREREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzN3d3dEREQzMzMiIiIiIiIREREiIiIREREiIiIiIiIiIiIREREiIiIREREiIiIREREREREiIiIiIiJVVVWIiIhmZmZmZmZmZmZVVVVVVVVERERERERVVVVERERVVVVERERERERERERVVVVVVVVERERmZmZVVVVVVVVVVVVVVVVERERERERERERERERERERERERVVVVVVVVVVVVVVVVERERERERVVVVERERVVVVVVVVVVVV3d3d3d3dmZmZVVVVVVVVERERERERERERERERERERERERVVVVERERERERVVVVERERERERERERERERVVVVERERERERVVVVVVVVmZmZVVVVVVVV3d3eqqqrMzMyIiIhVVVVVVVVVVVVmZmZ3d3eZmZlmZmZmZmZmZmZVVVV3d3d3d3dVVVUzMzNEREQzMzNVVVWZmZmZmZl3d3dERERVVVVmZmZEREQiIiIREREiIiIiIiIzMzMiIiIzMzMzMzMzMzNEREQzMzMzMzNERERERERERERERERVVVVEREREREQzMzNEREREREREREQzMzNERERERERERERVVVVVVVVEREQzMzNERERERERVVVVERERERERERERERERERERERERERERERERERERERERERERVVVVVVVVEREREREQzMzNEREREREREREQzMzMzMzMzMzNERERERERVVVVVVVVVVVVVVVVEREREREREREREREQzMzNEREREREQzMzNERERERERERERVVVVVVVVERERVVVVmZmZVVVVVVVVmZmZmZmZERERERERERERVVVVERERVVVVmZmZmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVV3d3d3d3dERERERERERERERERVVVVERERVVVVVVVVERERERERERERERERERERERERVVVVVVVVVVVVmZmZmZmZVVVVmZmZVVVVmZmZ3d3dmZmZmZmZmZmZVVVVVVVVERERVVVVmZmZVVVUzMzMiIiJERERVVVVVVVVERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVUzMzMzMzNVVVWZmZmIiIiIiIiIiIhERERERERmZmaZmZl3d3dVVVV3d3eZmZl3d3dVVVVERERVVVV3d3dmZmZEREQzMzMzMzNERERERERERERERERERERERERVVVVmZmZ3d3dmZmZmZmZmZmZVVVVERERERERmZmZ3d3d3d3d3d3dmZmZmZmZ3d3eIiIiIiIiZmZmqqqpmZmZVVVVVVVVVVVVVVVV3d3fMzMzu7u67u7uZmZnd3d3d3d27u7t3d3dVVVVVVVVmZmZmZmZ3d3dmZmZVVVVVVVVERERVVVVVVVV3d3d3d3dEREREREREREREREQzMzNEREQzMzMzMzMzMzNERERERERERERVVVVVVVVmZmZmZmZmZmZVVVVVVVVERERERERERERERERERERmZmaZmZm7u7vMzMyZmZm7u7vd3d3u7u7u7u7////////////////////////u7u7////////u7u7///////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzM3d3d3d3dzMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7zMzM3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7u7u7zMzMu7u7u7u7u7u7zMzMu7u7u7u7u7u7u7u7u7u7qqqqqqqqqqqqqqqqmZmZqqqqmZmZmZmZmZmZmZmZiIiIiIiIiIiId3d3iIiIiIiIiIiImZmZmZmZmZmZqqqqqqqqqqqqmZmZqqqqqqqqqqqqqqqqqqqqmZmZiIiImZmZqqqqmZmZmZmZmZmZiIiImZmZmZmZmZmZmZmZmZmZiIiIiIiIiIiId3d3d3d3iIiId3d3d3d3d3d3iIiIiIiIiIiIiIiId3d3d3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVZmZmZmZmVVVVZmZmZmZmZmZmVVVVREREVVVVVVVVVVVVVVVVd3d3iIiId3d3ZmZmZmZmd3d3ZmZmZmZmd3d3d3d3ZmZmd3d3iIiIiIiId3d3d3d3ZmZmVVVVVVVVd3d3d3d3ZmZmd3d3iIiId3d3d3d3ZmZmiIiIiIiId3d3d3d3iIiId3d3ZmZmZmZmVVVVZmZmiIiIZmZmZmZmVVVVVVVVVVVVVVVVd3d3d3d3ZmZmVVVVREREVVVVVVVVREREREREMzMzREREREREREREREREVVVViIiIu7u7u7u7u7u7mZmZqqqqqqqqqqqqd3d3d3d3mZmZiIiIzMzMzMzMzMzMu7u7zMzMzMzMu7u7zMzMzMzMu7u7u7u7qqqqmZmZd3d3mZmZu7u7zMzMu7u7qqqqqqqqu7u7zMzMzMzMu7u7qqqqqqqqqqqqqqqqmZmZd3d3d3d3d3d3iIiId3d3d3d3d3d3qqqqzMzMu7u7u7u7qqqqzMzMzMzMzMzMzMzMu7u7u7u7u7u7qqqqmZmZmZmZd3d3ZmZmiIiImZmZqqqqzMzMu7u7qqqqqqqqzMzMzMzMu7u7u7u7u7u7iIiIiIiIiIiIiIiId3d3d3d3d3d3VVVVd3d3iIiImZmZu7u7u7u7u7u7u7u7u7u7qqqqiIiIiIiImZmZqqqqqqqqu7u7qqqqmZmZmZmZd3d3VVVVZmZmmZmZmZmZmZmZqqqqmZmZiIiIiIiIiIiId3d3ZmZmZmZmZmZmVVVVZmZmZmZmVVVVd3d3iIiImZmZmZmZiIiImZmZqqqqqqqqmZmZiIiImZmZiIiId3d3d3d3d3d3d3d3d3d3ZmZmVVVVd3d3u7u7u7u7u7u7qqqqqqqqqqqqqqqqmZmZmZmZiIiId3d3iIiIiIiId3d3ZmZmVVVVVVVVd3d3qqqqzMzMu7u7qqqqqqqqiIiIiIiIiIiIiIiIiIiImZmZd3d3d3d3iIiIiIiId3d3iIiIiIiImZmZzMzMu7u7mZmZZmZmVVVVREREREREREREZmZmZmZmVVVVVVVVVVVVREREVVVVZmZmiIiImZmZmZmZqqqqqqqqmZmZd3d3iIiIiIiId3d3d3d3mZmZiIiId3d3d3d3ZmZmREREREREREREREREREREMzMzVVVVZmZmiIiImZmZmZmZiIiIiIiIqqqqzMzMqqqqmZmZVVVVVVVVVVVVVVVVZmZmVVVVVVVVd3d3iIiId3d3d3d3VVVVREREZmZmd3d3d3d3qqqqmZmZiIiIiIiIZmZmVVVVVVVVZmZmVVVVVVVVVVVVZmZmd3d3d3d3ZmZmVVVVZmZmZmZmVVVVZmZmZmZmd3d3iIiIiIiId3d3d3d3d3d3ZmZmREREREREREREMzMzREREVVVVVVVVVVVVZmZmZmZmREREVVVVVVVVVVVViIiIu7u7qqqqmZmZd3d3d3d3ZmZmREREVVVVREREREREREREREREVVVVREREREREREREREREMzMzIiIiREREiIiImZmZd3d3d3d3d3d3ZmZmZmZmZmZmZmZmVVVVVVVVZmZmZmZmVVVVVVVVREREREREREREREREVVVVREREVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVREREZmZmZmZmZmZmVVVVVVVVVVVVREREREREVVVVVVVVREREVVVVVVVVREREVVVVZmZmVVVVREREREREMzMzMzMzREREREREREREREREMzMzMzMzMzMzMzMzREREREREREREIiIiREREVVVVVVVVZmZmd3d3ZmZmZmZmZmZmVVVVVVVVREREREREMzMzREREVVVVVVVVREREREREREREMzMzREREREREREREREREREREVVVVZmZmVVVVVVVVZmZmVVVVVVVVREREVVVVVVVVVVVVREREREREREREMzMzMzMzREREMzMzMzMzREREMzMzREREMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiREREd3d3REREIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiERERIiIiREREZmZmZmZmVVVVZmZmVVVVREREREREVVVVREREVVVVREREVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVREREVVVVREREVVVVVVVVREREREREREREVVVVVVVVVVVVREREREREVVVVREREREREREREREREVVVVVVVVVVVVVVVVREREMzMzREREREREREREREREREREREREVVVVREREMzMzREREMzMzMzMzREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVViIiIzMzMqqqqd3d3d3d3ZmZmREREVVVVd3d3d3d3VVVVVVVVVVVVVVVVZmZmZmZmREREMzMzMzMzMzMzREREd3d3iIiId3d3ZmZmZmZmZmZmMzMzERERERERIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzREREVVVVREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVREREREREREREVVVVVVVVMzMzREREREREREREREREMzMzREREREREREREREREVVVVVVVVVVVVVVVVVVVVREREREREVVVVREREMzMzMzMzMzMzREREREREVVVVREREREREREREREREVVVVREREREREREREREREMzMzREREREREVVVVVVVVVVVVVVVVREREVVVVZmZmZmZmVVVVZmZmZmZmVVVVVVVVVVVVREREREREZmZmd3d3VVVVZmZmZmZmZmZmZmZmVVVVREREVVVVd3d3VVVVREREREREREREREREREREVVVVREREREREREREMzMzREREREREVVVVVVVVVVVVVVVVZmZmd3d3ZmZmZmZmVVVVVVVVZmZmd3d3ZmZmZmZmVVVVVVVVZmZmZmZmVVVVZmZmZmZmREREMzMzMzMzREREREREMzMzREREREREVVVVREREVVVVREREVVVVVVVVVVVVMzMzREREMzMzVVVVZmZmiIiId3d3d3d3ZmZmmZmZiIiIVVVVREREREREZmZmiIiId3d3REREREREVVVVZmZmVVVVREREREREREREREREVVVVVVVVVVVVREREVVVVZmZmZmZmd3d3d3d3d3d3VVVVREREVVVVZmZmd3d3d3d3ZmZmZmZmZmZmd3d3mZmZqqqqu7u7qqqqZmZmVVVVREREVVVVVVVVd3d3zMzM7u7uzMzMqqqqzMzMzMzMiIiId3d3VVVVVVVVd3d3iIiIiIiIiIiId3d3VVVVREREREREVVVVVVVVZmZmREREREREREREREREREREMzMzMzMzREREREREREREMzMzREREREREVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVREREREREREREZmZmiIiIqqqqqqqqmZmZqqqqzMzM3d3d3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7t3d3czMzMzMzMzMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzLu7u7u7u7u7u7u7u8zMzMzMzMzMzMzMzMzMzLu7u8zMzLu7u7u7u7u7u7u7u6qqqru7u6qqqqqqqru7u7u7u7u7u7u7u7u7u6qqqpmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiJmZmYiIiIiIiIiIiJmZmYiIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiHd3d3d3d4iIiHd3d4iIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiHd3d4iIiJmZmZmZmYiIiHd3d3d3d3d3d4iIiHd3d4iIiIiIiHd3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVURERERERERERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERERERFVVVXd3d3d3d2ZmZmZmZnd3d2ZmZmZmZmZmZlVVVWZmZmZmZnd3d4iIiHd3d3d3d2ZmZlVVVVVVVWZmZnd3d2ZmZmZmZoiIiIiIiHd3d3d3d3d3d4iIiIiIiIiIiHd3d3d3d3d3d3d3d2ZmZnd3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVWZmZmZmZlVVVWZmZlVVVURERFVVVURERERERERERERERFVVVTMzM1VVVXd3d5mZmbu7u8zMzMzMzMzMzLu7u7u7u7u7u4iIiJmZmZmZmaqqqszMzMzMzLu7u7u7u93d3czMzLu7u6qqqszMzLu7u6qqqqqqqoiIiIiIiIiIiLu7u8zMzLu7u6qqqru7u7u7u7u7u7u7u7u7u5mZmZmZmaqqqqqqqoiIiHd3d3d3d3d3d4iIiGZmZnd3d4iIiKqqqszMzLu7u5mZmaqqqru7u93d3czMzMzMzLu7u7u7u8zMzLu7u7u7u5mZmXd3d3d3d4iIiJmZmZmZmbu7u8zMzKqqqqqqqru7u7u7u7u7u7u7u6qqqoiIiJmZmZmZmYiIiIiIiJmZmYiIiGZmZmZmZpmZmaqqqszMzMzMzMzMzLu7u6qqqqqqqqqqqpmZmZmZmZmZmZmZmaqqqru7u6qqqpmZmYiIiGZmZmZmZpmZmZmZmZmZmZmZmXd3d4iIiHd3d2ZmZmZmZnd3d3d3d2ZmZlVVVXd3d4iIiGZmZmZmZoiIiJmZmZmZmaqqqpmZmaqqqqqqqpmZmZmZmYiIiHd3d3d3d3d3d3d3d3d3d3d3d1VVVVVVVWZmZqqqqru7u7u7u6qqqqqqqqqqqqqqqqqqqoiIiIiIiIiIiIiIiIiIiGZmZmZmZmZmZmZmZnd3d4iIiKqqqru7u6qqqoiIiIiIiKqqqpmZmYiIiIiIiIiIiHd3d3d3d5mZmYiIiIiIiIiIiGZmZoiIiLu7u6qqqoiIiGZmZlVVVURERERERFVVVVVVVWZmZmZmZkRERFVVVVVVVWZmZnd3d4iIiJmZmZmZmZmZmbu7u5mZmXd3d4iIiIiIiGZmZnd3d4iIiHd3d4iIiHd3d2ZmZkRERERERERERERERDMzM0RERERERFVVVWZmZoiIiJmZmYiIiIiIiLu7u7u7u6qqqnd3d1VVVVVVVVVVVWZmZmZmZmZmZkRERGZmZoiIiHd3d4iIiGZmZkRERFVVVVVVVXd3d6qqqpmZmZmZmYiIiHd3d1VVVVVVVWZmZlVVVVVVVVVVVVVVVWZmZnd3d1VVVVVVVWZmZlVVVVVVVWZmZoiIiJmZmYiIiIiIiHd3d3d3d3d3d3d3d1VVVVVVVVVVVURERERERERERFVVVVVVVVVVVVVVVVVVVURERFVVVVVVVYiIiJmZmZmZmYiIiHd3d2ZmZmZmZmZmZlVVVVVVVVVVVWZmZlVVVURERERERERERERERDMzMzMzMyIiIkRERHd3d4iIiHd3d3d3d3d3d3d3d2ZmZlVVVVVVVVVVVWZmZlVVVWZmZmZmZlVVVVVVVVVVVVVVVURERFVVVURERFVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVURERGZmZmZmZmZmZlVVVURERGZmZlVVVVVVVWZmZkRERERERERERFVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERERERERERERERDMzM0RERERERERERDMzMzMzMzMzM0RERERERGZmZmZmZmZmZmZmZlVVVVVVVVVVVURERERERERERERERFVVVVVVVVVVVURERERERERERERERERERERERERERDMzM1VVVXd3d2ZmZkRERFVVVVVVVVVVVVVVVVVVVURERFVVVVVVVURERERERERERERERERERERERDMzM0RERERERERERDMzMzMzMyIiIiIiIjMzMzMzMyIiIiIiIjMzM2ZmZjMzMyIiIiIiIiIiIhERESIiIhERESIiIhERESIiIhERERERESIiIiIiIiIiIiIiIiIiIiIiIjMzM1VVVWZmZmZmZmZmZlVVVVVVVVVVVURERERERERERFVVVVVVVVVVVURERFVVVVVVVWZmZlVVVURERERERFVVVURERFVVVVVVVWZmZlVVVVVVVURERERERFVVVURERERERERERERERERERERERERERERERERERERERERERERERERERDMzM0RERERERDMzM0RERERERFVVVURERERERDMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVVVVVWZmZlVVVVVVVVVVVWZmZpmZmczMzIiIiHd3d5mZmXd3d1VVVVVVVXd3d2ZmZlVVVVVVVURERFVVVWZmZlVVVURERDMzMzMzMzMzM0RERHd3d5mZmYiIiGZmZmZmZlVVVTMzMyIiIhERERERESIiIhERESIiIiIiIjMzMzMzMzMzM0RERERERDMzMzMzM0RERERERERERFVVVURERERERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVTMzM0RERERERERERDMzM0RERERERERERERERERERERERFVVVVVVVVVVVVVVVURERFVVVWZmZlVVVTMzMzMzM0RERERERFVVVURERFVVVVVVVURERERERERERFVVVURERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVWZmZmZmZkRERERERGZmZkRERERERIiIiIiIiGZmZnd3d3d3d3d3d2ZmZlVVVVVVVVVVVWZmZmZmZkRERERERERERERERFVVVURERERERERERERERDMzMzMzM0RERGZmZlVVVURERFVVVXd3d2ZmZnd3d1VVVWZmZmZmZlVVVYiIiHd3d2ZmZlVVVXd3d4iIiHd3d2ZmZlVVVVVVVVVVVTMzMzMzMzMzMzMzM0RERERERERERERERFVVVURERERERFVVVVVVVVVVVURERDMzMzMzM0RERERERFVVVWZmZlVVVVVVVWZmZmZmZnd3d4iIiHd3d1VVVXd3d3d3d1VVVURERERERERERERERDMzM0RERERERERERERERERERFVVVVVVVVVVVWZmZnd3d2ZmZmZmZlVVVURERERERGZmZnd3d3d3d3d3d3d3d2ZmZmZmZnd3d3d3d5mZmaqqqpmZmXd3d1VVVURERERERGZmZmZmZqqqqu7u7ru7u6qqqt3d3d3d3ZmZmYiIiHd3d2ZmZoiIiIiIiIiIiIiIiHd3d3d3d2ZmZlVVVVVVVURERFVVVVVVVURERERERERERERERERERERERDMzM0RERDMzM0RERERERERERERERERERFVVVVVVVVVVVURERERERFVVVVVVVURERERERERERHd3d6qqqpmZmYiIiKqqqszMzMzMzO7u7t3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3u7u7d3d3u7u7d3d3u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3d3d3d3d3MzMzMzMzMzMzMzMy7u7u7u7u7u7vMzMy7u7u7u7vMzMy7u7u7u7u7u7u7u7u7u7uqqqq7u7uqqqqqqqqqqqqqqqqqqqqZmZmIiIiIiIh3d3eIiIiIiIh3d3eIiIiIiIiIiIiIiIiZmZmIiIiIiIiIiIiZmZmZmZmZmZmZmZmIiIiZmZmZmZmZmZmIiIiZmZmIiIiIiIiIiIiIiIiIiIh3d3eIiIh3d3dmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3eIiIiIiIh3d3d3d3eIiIh3d3eIiIiZmZmIiIh3d3d3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZVVVVVVVVVVVVVVVVERERVVVVERERERERVVVVmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3dVVVVERERmZmZmZmZmZmZmZmaIiIh3d3dmZmZ3d3eIiIiZmZmqqqqIiIh3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3d3d3eIiIh3d3dmZmZVVVVVVVVVVVVVVVV3d3dmZmZmZmZEREREREREREREREQzMzNEREQzMzNmZmZ3d3eZmZm7u7vd3d3MzMzMzMzMzMy7u7uqqqqIiIiqqqq7u7vMzMzMzMzMzMzMzMzd3d3d3d3MzMy7u7uqqqq7u7u7u7uqqqqZmZmZmZl3d3dmZmaZmZm7u7u7u7uqqqqqqqq7u7uqqqq7u7u7u7uqqqqZmZmqqqqZmZmIiIh3d3eIiIh3d3d3d3dmZmZ3d3eZmZm7u7vMzMzMzMyqqqq7u7u7u7vMzMzMzMzMzMzMzMyqqqqqqqq7u7uqqqqqqqqIiIiIiIiZmZmIiIiZmZm7u7vMzMzMzMy7u7u7u7vMzMy7u7uqqqqZmZmqqqq7u7uqqqqZmZmqqqqqqqqZmZl3d3dmZmZ3d3eZmZnMzMzMzMzd3d27u7uqqqqqqqqqqqqqqqq7u7uZmZmIiIiZmZmqqqq7u7uqqqqqqqqIiIhmZmaIiIiZmZmqqqqZmZmqqqqZmZl3d3eIiIh3d3d3d3dmZmZmZmZVVVVVVVV3d3dmZmZVVVVmZmZ3d3eIiIiZmZmZmZmZmZmqqqqZmZmIiIiIiIiIiIh3d3dmZmZ3d3d3d3dmZmZmZmZ3d3dmZmaZmZmqqqq7u7uqqqqqqqqqqqqZmZmZmZmZmZmIiIiZmZl3d3dmZmZmZmZmZmZ3d3dmZmZ3d3eIiIiZmZmqqqqZmZmZmZmqqqqqqqqIiIiqqqqZmZmIiIiIiIiIiIiZmZmIiIiIiIh3d3dVVVVmZmaZmZmZmZlmZmZmZmZVVVVVVVVVVVVERERVVVVmZmZVVVVVVVVVVVVmZmZ3d3d3d3eIiIiZmZmqqqqZmZmqqqq7u7uZmZmIiIh3d3d3d3d3d3d3d3eIiIiZmZmIiIhVVVVERERERERVVVVERERERERERERERERVVVVmZmZmZmZmZmZmZmaZmZm7u7u7u7uZmZlmZmZVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVV3d3eIiIiIiIh3d3dmZmZERERmZmaZmZmZmZmZmZl3d3d3d3dmZmZmZmZmZmZ3d3dmZmZVVVVERERVVVVmZmZ3d3dmZmZmZmZmZmZVVVVVVVV3d3d3d3eZmZmZmZmZmZmIiIh3d3d3d3dmZmZVVVVmZmZmZmZVVVVERERERERERERVVVVmZmZVVVVERERVVVVVVVVmZmaZmZmZmZmZmZmZmZl3d3d3d3d3d3dmZmZmZmZmZmZVVVVVVVVVVVVVVVVEREREREREREREREREREQzMzNERER3d3eIiIh3d3d3d3dmZmZ3d3dmZmZmZmZVVVVmZmZVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZVVVV3d3dmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERERERVVVVVVVVVVVVVVVVEREREREREREQzMzMzMzNERERVVVVEREREREREREREREREREREREREREREREREREQzMzMzMzNERERVVVVmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVmZmZVVVVmZmZmZmZERERVVVVEREREREQzMzNERERmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVmZmZVVVVEREQzMzMzMzMiIiIzMzMzMzMiIiIiIiIiIiIzMzNEREQzMzMiIiIREREiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiJERERmZmZmZmZmZmZVVVVmZmZVVVVERERVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERVVVVVVVVERERVVVVVVVVERERVVVVVVVVVVVVEREREREREREREREQzMzMzMzNEREQzMzNEREQzMzNEREREREQzMzNEREQzMzMzMzNEREREREREREREREREREREREQzMzMzMzMzMzMzMzNEREQzMzNVVVVVVVVVVVVVVVVVVVVVVVVVVVWIiIiqqqqZmZlmZmZ3d3eqqqqZmZlERERmZmZ3d3dVVVVERERERERERERERERVVVVEREQzMzMzMzMzMzMzMzNERER3d3eqqqqZmZlmZmZVVVVmZmZEREQiIiIREREREREiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVERERERERERERERERERERVVVVERERVVVVERERVVVVmZmZmZmZVVVVVVVVERERVVVVVVVUzMzNEREREREREREREREQzMzNEREQzMzNERERERERERERERERVVVVERERVVVVVVVVVVVVmZmZmZmZERERERERERERERERERERVVVVVVVVVVVVmZmZVVVVVVVVERERVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmIiIiqqqqqqqp3d3d3d3dmZmZVVVVERERVVVVmZmZERERERERERERVVVVEREREREQzMzMzMzMzMzMzMzMzMzNERERmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmaIiIiIiIiIiIhmZmZ3d3eZmZmqqqp3d3dmZmZVVVVmZmZEREQzMzMzMzMzMzNERERERERVVVVERERERERERERVVVVERERVVVVEREREREREREREREQzMzNEREREREREREQzMzMzMzNERERmZmaZmZm7u7uZmZl3d3dmZmZmZmZmZmZVVVVEREQzMzMzMzMzMzNERERERERVVVVVVVVERERVVVVmZmZmZmZmZmZmZmZmZmZERERERERERERVVVV3d3d3d3d3d3d3d3dmZmZVVVVmZmZmZmZmZmaIiIh3d3dmZmZmZmZVVVVERER3d3eZmZl3d3eIiIi7u7u7u7u7u7vd3d3u7u67u7vMzMy7u7uIiIh3d3eqqqq7u7uZmZlmZmZmZmZmZmZVVVVERERVVVVERERVVVVmZmZVVVVEREREREREREREREREREREREREREREREQzMzNERERERERERERVVVVVVVVEREREREQzMzNERERmZmZVVVVERERERER3d3eZmZl3d3dmZmaZmZm7u7vd3d3d3d3d3d3d3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////7u7u7u7u3d3d3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3dzMzMzMzMzMzMzMzM3d3d3d3d3d3d3d3d7u7u7u7u7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3d3d3dzMzM3d3dzMzMzMzM3d3dzMzM3d3d3d3dzMzMzMzMzMzMzMzMzMzMu7u7zMzMzMzMzMzMzMzMu7u7zMzMu7u7u7u7qqqqqqqqmZmZqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqmZmZmZmZmZmZmZmZqqqqmZmZiIiIiIiIiIiId3d3d3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiId3d3iIiId3d3iIiId3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3d3d3iIiIiIiId3d3d3d3d3d3iIiId3d3iIiId3d3d3d3d3d3d3d3d3d3ZmZmZmZmd3d3ZmZmZmZmZmZmZmZmd3d3iIiId3d3ZmZmd3d3d3d3d3d3d3d3d3d3ZmZmd3d3iIiId3d3VVVVVVVVd3d3ZmZmZmZmd3d3ZmZmZmZmd3d3d3d3iIiIqqqqiIiId3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiId3d3iIiId3d3ZmZmZmZmZmZmVVVVVVVVd3d3ZmZmVVVVREREREREREREMzMzREREREREMzMzVVVVd3d3mZmZzMzMu7u7zMzMu7u7qqqqqqqqiIiIiIiIu7u7zMzMzMzMu7u7zMzM3d3d3d3d3d3d3d3dzMzMqqqqqqqqu7u7u7u7mZmZiIiIZmZmVVVVd3d3qqqqzMzMqqqqqqqqzMzMu7u7u7u7u7u7qqqqiIiImZmZmZmZiIiIiIiId3d3VVVVVVVVZmZmd3d3mZmZqqqqzMzMzMzMzMzMu7u7u7u7u7u7zMzMzMzMu7u7qqqqmZmZmZmZqqqqmZmZmZmZmZmZqqqqmZmZiIiIu7u7zMzM3d3du7u7u7u7u7u7u7u7u7u7qqqqzMzMu7u7qqqqqqqqmZmZqqqqiIiId3d3d3d3ZmZmZmZmmZmZu7u7u7u7u7u7u7u7qqqqqqqqmZmZqqqqmZmZiIiImZmZqqqqqqqqmZmZmZmZiIiId3d3d3d3qqqqu7u7qqqqu7u7qqqqmZmZiIiIiIiIVVVVVVVVZmZmZmZmREREVVVVZmZmd3d3d3d3d3d3iIiIiIiIiIiIqqqqqqqqmZmZiIiIiIiIiIiId3d3d3d3d3d3ZmZmVVVVZmZmd3d3d3d3d3d3qqqqu7u7u7u7qqqqqqqqmZmZiIiIiIiImZmZmZmZd3d3VVVVZmZmiIiIZmZmZmZmd3d3iIiImZmZqqqqqqqqmZmZmZmZiIiImZmZmZmZmZmZmZmZmZmZd3d3mZmZiIiIiIiId3d3ZmZmd3d3iIiIiIiId3d3iIiId3d3VVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmd3d3iIiImZmZmZmZmZmZmZmZmZmZmZmZu7u7mZmZiIiIiIiId3d3d3d3d3d3iIiIiIiIZmZmVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmVVVVZmZmmZmZu7u7qqqqiIiIZmZmVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmiIiId3d3iIiIiIiId3d3ZmZmd3d3mZmZqqqqmZmZd3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmVVVVVVVVd3d3d3d3ZmZmZmZmZmZmZmZmVVVVd3d3iIiIiIiIiIiImZmZmZmZd3d3ZmZmZmZmVVVVVVVVVVVVVVVVREREREREREREZmZmVVVVVVVVREREREREVVVVZmZmmZmZqqqqmZmZiIiIiIiIZmZmd3d3ZmZmZmZmZmZmVVVVREREVVVVZmZmZmZmVVVVVVVVVVVVVVVVMzMzMzMzZmZmiIiIiIiId3d3ZmZmVVVVZmZmZmZmZmZmVVVVVVVVZmZmZmZmd3d3ZmZmZmZmZmZmZmZmd3d3d3d3ZmZmREREZmZmZmZmVVVVd3d3ZmZmVVVVVVVVZmZmZmZmVVVVVVVVZmZmZmZmZmZmVVVVZmZmVVVVZmZmZmZmVVVVVVVVREREMzMzVVVVVVVVZmZmZmZmVVVVVVVVREREREREREREREREREREREREREREVVVVZmZmVVVVREREREREVVVVVVVVREREREREREREVVVVZmZmZmZmREREZmZmZmZmVVVVVVVVVVVVVVVVVVVVREREREREVVVVREREVVVVVVVVVVVVd3d3VVVVVVVVVVVVREREMzMzVVVVZmZmVVVVREREZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVREREVVVVVVVVREREVVVVZmZmd3d3ZmZmVVVVREREREREREREMzMzMzMzMzMzMzMzIiIiIiIiMzMzREREMzMzIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiREREZmZmZmZmZmZmVVVVVVVVZmZmVVVVVVVVREREVVVVREREREREVVVVREREVVVVREREREREREREREREVVVVVVVVREREVVVVREREVVVVREREVVVVREREVVVVVVVVVVVVREREREREMzMzREREMzMzREREMzMzREREREREREREREREREREREREREREMzMzMzMzREREREREREREREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVViIiIu7u7iIiIVVVVZmZmd3d3ZmZmREREZmZmZmZmVVVVREREMzMzMzMzMzMzMzMzREREMzMzIiIiMzMzMzMzMzMzVVVVmZmZmZmZZmZmd3d3d3d3REREIiIiIiIiIiIiERERIiIiIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzREREMzMzREREREREMzMzMzMzREREREREREREREREREREVVVVREREVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREREREMzMzREREREREREREREREMzMzREREREREREREREREREREREREVVVVVVVVVVVVVVVVd3d3ZmZmREREREREREREREREVVVVVVVVVVVVZmZmZmZmZmZmVVVVREREREREVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVd3d3mZmZiIiIiIiIzMzMzMzMiIiId3d3mZmZZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREMzMzREREMzMzMzMzMzMzMzMzREREVVVVZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVZmZmiIiImZmZiIiImZmZmZmZqqqqmZmZd3d3VVVVVVVVZmZmVVVVMzMzIiIiREREMzMzVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREREREREREREREREREMzMzREREMzMzREREd3d3mZmZqqqqmZmZd3d3ZmZmVVVVZmZmZmZmREREREREMzMzMzMzREREVVVVVVVVZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmVVVVREREREREZmZmd3d3ZmZmd3d3d3d3d3d3ZmZmVVVVZmZmZmZmd3d3d3d3REREREREZmZmZmZmVVVVZmZmqqqqmZmZiIiImZmZu7u7zMzM3d3d7u7u3d3d7u7u7u7uqqqqZmZmmZmZu7u7mZmZZmZmZmZmREREVVVVREREREREVVVVVVVVZmZmVVVVVVVVREREREREVVVVREREREREREREREREREREMzMzREREREREREREREREREREMzMzMzMzMzMzREREVVVVVVVVVVVVd3d3iIiIVVVVREREd3d3qqqqzMzM3d3d3d3d3d3d3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7t3d3d3d3d3d3e7u7u7u7t3d3e7u7t3d3d3d3d3d3czMzN3d3czMzMzMzMzMzMzMzMzMzLu7u8zMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u8zMzLu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqqqqqqqqqqqqqqqqqru7u7u7u6qqqqqqqqqqqqqqqqqqqru7u6qqqpmZmaqqqqqqqpmZmaqqqqqqqqqqqpmZmaqqqqqqqpmZmZmZmaqqqpmZmYiIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiIiIiIiIiIiIiJmZmZmZmZmZmZmZmYiIiIiIiIiIiIiIiHd3d4iIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiHd3d4iIiIiIiHd3d4iIiHd3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d2ZmZnd3d2ZmZmZmZmZmZnd3d3d3d3d3d2ZmZlVVVWZmZnd3d2ZmZnd3d4iIiHd3d2ZmZmZmZmZmZoiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d4iIiIiIiHd3d5mZmYiIiHd3d2ZmZmZmZmZmZmZmZmZmZnd3d1VVVVVVVURERDMzMzMzM0RERFVVVURERERERGZmZoiIiKqqqszMzLu7u6qqqru7u6qqqru7u4iIiJmZmczMzN3d3bu7u6qqqszMzN3d3e7u7u7u7t3d3czMzKqqqru7u8zMzKqqqoiIiIiIiGZmZlVVVXd3d6qqqszMzLu7u6qqqru7u8zMzLu7u5mZmYiIiJmZmYiIiIiIiIiIiIiIiGZmZlVVVVVVVXd3d4iIiIiIiKqqqszMzMzMzLu7u6qqqqqqqru7u8zMzMzMzLu7u6qqqoiIiJmZmZmZmYiIiIiIiIiIiJmZmZmZmYiIiJmZmczMzN3d3czMzLu7u7u7u6qqqru7u7u7u7u7u6qqqqqqqpmZmZmZmYiIiIiIiIiIiIiIiHd3d2ZmZnd3d7u7u8zMzLu7u7u7u7u7u6qqqpmZmZmZmYiIiIiIiIiIiLu7u5mZmXd3d4iIiJmZmYiIiHd3d5mZmbu7u7u7u6qqqpmZmXd3d3d3d2ZmZlVVVWZmZmZmZmZmZlVVVURERGZmZoiIiJmZmYiIiIiIiIiIiJmZmaqqqqqqqpmZmYiIiHd3d3d3d4iIiIiIiFVVVWZmZmZmZmZmZmZmZmZmZoiIiKqqqru7u7u7u6qqqqqqqoiIiIiIiJmZmYiIiIiIiGZmZnd3d3d3d3d3d2ZmZnd3d3d3d4iIiIiIiJmZmbu7u7u7u5mZmZmZmZmZmYiIiJmZmaqqqpmZmXd3d4iIiJmZmZmZmYiIiHd3d5mZmaqqqoiIiGZmZnd3d4iIiGZmZlVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d4iIiIiIiKqqqpmZmZmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiHd3d3d3d3d3d4iIiIiIiFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZoiIiKqqqqqqqqqqqoiIiHd3d2ZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d4iIiIiIiHd3d3d3d2ZmZmZmZnd3d4iIiJmZmZmZmYiIiHd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZlVVVWZmZnd3d5mZmYiIiIiIiIiIiIiIiGZmZmZmZnd3d2ZmZlVVVWZmZmZmZlVVVVVVVVVVVWZmZlVVVVVVVURERERERDMzM1VVVZmZmaqqqoiIiHd3d4iIiHd3d2ZmZmZmZmZmZlVVVWZmZlVVVVVVVWZmZmZmZlVVVWZmZmZmZlVVVURERDMzM2ZmZoiIiIiIiHd3d2ZmZmZmZlVVVWZmZmZmZlVVVWZmZmZmZmZmZnd3d2ZmZmZmZnd3d4iIiIiIiHd3d0RERERERGZmZmZmZlVVVWZmZmZmZlVVVWZmZlVVVVVVVWZmZmZmZmZmZlVVVWZmZmZmZlVVVWZmZlVVVVVVVWZmZlVVVURERERERFVVVVVVVVVVVWZmZlVVVURERERERFVVVVVVVURERFVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVURERERERERERGZmZnd3d2ZmZlVVVWZmZlVVVVVVVVVVVVVVVURERFVVVURERERERERERFVVVWZmZlVVVWZmZmZmZlVVVVVVVVVVVURERERERFVVVWZmZlVVVVVVVWZmZlVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVURERERERFVVVWZmZnd3d2ZmZlVVVVVVVVVVVURERDMzMzMzMzMzMzMzMyIiIiIiIkRERFVVVURERCIiIjMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIkRERFVVVXd3d2ZmZlVVVWZmZlVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERERERFVVVVVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERDMzMzMzM0RERERERERERERERERERERERERERERERERERDMzMzMzM0RERERERDMzM0RERDMzM0RERERERERERERERDMzM0RERDMzM0RERFVVVVVVVVVVVWZmZmZmZnd3d5mZmaqqqnd3d0RERFVVVVVVVURERFVVVWZmZlVVVURERDMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzM1VVVZmZmZmZmXd3d3d3d2ZmZkRERDMzMxERERERERERESIiIiIiIjMzMyIiIjMzMyIiIiIiIjMzMzMzMzMzMzMzM0RERDMzM0RERERERERERERERFVVVVVVVURERFVVVURERFVVVVVVVWZmZlVVVVVVVURERFVVVURERDMzM0RERERERERERDMzM0RERERERERERERERERERDMzM0RERERERFVVVWZmZlVVVVVVVXd3d1VVVVVVVURERFVVVURERERERFVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVURERFVVVVVVVWZmZnd3d3d3d2ZmZnd3d4iIiIiIiJmZmczMzMzMzHd3d4iIiKqqqmZmZlVVVURERFVVVVVVVVVVVURERERERERERERERDMzMzMzMzMzM0RERDMzM0RERFVVVWZmZmZmZlVVVURERFVVVVVVVVVVVVVVVWZmZlVVVWZmZnd3d4iIiJmZmaqqqqqqqqqqqqqqqnd3d2ZmZlVVVWZmZlVVVURERDMzMzMzMzMzM0RERFVVVVVVVURERFVVVURERERERERERERERERERERERERERERERERERERERERERERERERERFVVVXd3d4iIiJmZmXd3d2ZmZmZmZlVVVVVVVVVVVURERERERERERERERFVVVWZmZmZmZmZmZmZmZnd3d2ZmZmZmZlVVVURERERERFVVVWZmZnd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZoiIiGZmZkRERFVVVWZmZnd3d3d3d3d3d3d3d4iIiHd3d4iIiJmZmaqqqszMzN3d3d3d3e7u7t3d3aqqqnd3d3d3d6qqqru7u6qqqmZmZkRERFVVVURERERERERERFVVVVVVVVVVVVVVVURERFVVVURERERERFVVVURERERERERERERERERERERERERERDMzMzMzMzMzM0RERDMzM0RERFVVVVVVVVVVVXd3d2ZmZkRERERERGZmZoiIiLu7u93d3d3d3d3d3czMzN3d3e7u7v///////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3MzMzMzMzMzMzMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMy7u7vMzMyqqqq7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7uqqqqqqqq7u7uqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqZmZmZmZmZmZmIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZmIiIiIiIiIiIiIiIh3d3eIiIh3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3dmZmZ3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVmZmZVVVVVVVVVVVVmZmZmZmZ3d3dmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3eIiIh3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3eIiIiIiIiIiIh3d3d3d3dmZmZ3d3d3d3eIiIiZmZmIiIh3d3dmZmZ3d3d3d3dmZmZmZmZmZmZ3d3dVVVVEREREREREREQzMzNERERVVVVERERmZmaIiIiZmZm7u7u7u7u7u7uZmZmqqqrMzMy7u7uqqqqqqqqqqqq7u7u7u7u7u7vMzMzd3d3d3d3d3d3d3d27u7u7u7u7u7u7u7uqqqqIiIiIiIh3d3dVVVV3d3eqqqq7u7uqqqqqqqq7u7u7u7u7u7uIiIh3d3eIiIiZmZmIiIiZmZmZmZlmZmZVVVV3d3eIiIiZmZmIiIiIiIi7u7vMzMy7u7uqqqq7u7u7u7u7u7vMzMy7u7uqqqqIiIiIiIiZmZmIiIh3d3eIiIiZmZmZmZmIiIh3d3eqqqrd3d3MzMzMzMy7u7uqqqqqqqqqqqqqqqqqqqqqqqqZmZmZmZmIiIiIiIiZmZmqqqq7u7uIiIhmZmZ3d3e7u7vd3d3MzMy7u7u7u7u7u7uZmZmIiIh3d3eZmZmZmZmIiIh3d3eIiIiZmZmZmZl3d3eZmZm7u7uqqqqqqqqIiIh3d3d3d3dmZmZVVVVVVVV3d3dmZmZVVVVVVVVmZmaIiIiZmZmZmZmZmZmIiIiqqqq7u7uqqqqqqqqIiIiIiIiIiIiIiIhmZmZmZmZ3d3dmZmZmZmZ3d3d3d3d3d3eZmZm7u7vMzMzMzMyqqqqZmZmZmZmZmZmZmZl3d3d3d3d3d3eIiIh3d3eIiIh3d3d3d3d3d3eIiIiIiIiZmZm7u7u7u7uZmZmqqqqZmZmqqqqZmZl3d3d3d3eIiIiIiIiZmZmIiIiIiIiqqqqqqqp3d3dmZmZ3d3eIiIiIiIh3d3dmZmZVVVVVVVVVVVVmZmZmZmZ3d3eIiIiIiIiZmZmZmZmZmZmZmZmZmZmqqqqZmZmIiIiIiIh3d3eIiIiIiIh3d3eIiIh3d3dVVVVERERVVVVVVVVVVVVERERVVVVVVVVmZmZ3d3dmZmaIiIiZmZm7u7uqqqqIiIh3d3eIiIiIiIh3d3d3d3dmZmZmZmZ3d3d3d3eIiIiZmZmIiIh3d3d3d3dmZmZmZmZ3d3eIiIiqqqqZmZmIiIiIiIiIiIh3d3d3d3d3d3d3d3dmZmZ3d3eIiIh3d3d3d3dmZmZmZmZ3d3dVVVVVVVV3d3eZmZmZmZmZmZmIiIiIiIh3d3eIiIhmZmZVVVVmZmZ3d3dmZmZVVVVmZmZmZmZmZmZmZmZVVVVEREQzMzNERERERESIiIiZmZmIiIh3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZVVVVmZmZVVVUzMzMzMzNVVVWIiIiZmZl3d3d3d3dmZmZ3d3dmZmZ3d3d3d3dmZmZmZmZmZmZ3d3d3d3d3dwD//wAAd4iIiHd3d2ZmZmZmZkRERERERFVVVWZmZlVVVWZmZmZmZlVVVWZmZmZmZlVVVWZmZmZmZmZmZlVVVWZmZlVVVVVVVVVVVVVVVWZmZmZmZlVVVURERERERFVVVWZmZlVVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERERERDMzM0RERGZmZnd3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVURERFVVVURERFVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVWZmZlVVVURERDMzM1VVVWZmZmZmZlVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVXd3d2ZmZnd3d2ZmZmZmZlVVVURERDMzMzMzMzMzMzMzMyIiIiIiIkRERFVVVURERCIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIjMzMzMzM1VVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVURERERERERERERERDMzM0RERERERERERFVVVVVVVVVVVWZmZlVVVURERERERFVVVVVVVWZmZlVVVVVVVVVVVWZmZmZmZkRERERERDMzM0RERERERERERDMzM0RERDMzMzMzM0RERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVURERERERERERDMzMzMzM0RERFVVVVVVVWZmZlVVVXd3d5mZmaqqqoiIiGZmZlVVVURERFVVVWZmZmZmZlVVVVVVVTMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMyIiIjMzMzMzM0RERERERHd3d5mZmZmZmZmZmXd3d0RERDMzMyIiIiIiIhERESIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERFVVVURERFVVVVVVVURERFVVVVVVVWZmZlVVVVVVVURERERERERERERERDMzM0RERDMzM0RERERERDMzM0RERDMzM0RERERERFVVVVVVVWZmZlVVVVVVVVVVVWZmZlVVVVVVVURERERERERERFVVVVVVVVVVVVVVVVVVVWZmZlVVVURERFVVVVVVVVVVVURERFVVVWZmZnd3d3d3d2ZmZlVVVVVVVVVVVWZmZlVVVVVVVURERFVVVWZmZnd3d2ZmZnd3d4iIiHd3d5mZmaqqqszMzMzMzGZmZnd3d5mZmWZmZlVVVVVVVVVVVVVVVVVVVURERERERERERERERDMzM0RERDMzM0RERERERERERERERGZmZmZmZkRERERERERERERERFVVVVVVVVVVVVVVVWZmZmZmZmZmZoiIiKqqqru7u8zMzLu7u5mZmXd3d1VVVVVVVVVVVVVVVVVVVTMzMzMzMzMzM0RERERERFVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERERERFVVVURERERERGZmZnd3d3d3d3d3d3d3d2ZmZkRERERERERERFVVVVVVVURERERERFVVVWZmZmZmZmZmZnd3d3d3d2ZmZlVVVURERFVVVVVVVWZmZmZmZmZmZnd3d2ZmZmZmZlVVVWZmZmZmZlVVVWZmZoiIiGZmZlVVVVVVVWZmZoiIiIiIiIiIiHd3d2ZmZlVVVWZmZoiIiKqqqszMzN3d3d3d3e7u7u7u7szMzHd3d2ZmZqqqqt3d3aqqqoiIiGZmZkRERERERDMzM0RERFVVVVVVVVVVVURERFVVVVVVVURERFVVVURERFVVVURERERERERERERERERERERERDMzMzMzMzMzMzMzM0RERDMzM0RERERERGZmZmZmZlVVVTMzM0RERERERGZmZpmZmczMzO7u7t3d3d3d3czMzMzMzO7u7v///////+7u7v///////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7d3d3d3d3u7u7u7u7d3d3u7u7u7u7u7u7u7u7d3d3u7u7d3d3u7u7d3d3u7u7d3d3u7u7d3d3u7u7d3d3u7u7d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7uqqqq7u7u7u7uqqqqZmZmZmZmZmZmZmZmIiIiZmZmZmZmIiIiIiIiIiIh3d3eIiIiIiIh3d3dmZmZ3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVEREREREREREREREREREREREREREQzMzNEREREREQzMzNERERERERVVVVVVVVVVVVERERVVVVVVVVVVVVERERVVVVERERERERERERERERERERERERERERERERERERERERERERERERERERERERVVVVEREREREQzMzNEREQzMzNEREQzMzMzMzMzMzNEREQzMzNERERERERERERVVVVERERVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVV3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZ3d3eIiIh3d3d3d3d3d3dmZmZ3d3eIiIiIiIiIiIh3d3dmZmZ3d3d3d3dmZmZVVVVmZmZ3d3d3d3dmZmZmZmZVVVVERERVVVVVVVVmZmaZmZmZmZmIiIiZmZm7u7u7u7u7u7u7u7uqqqqZmZmZmZmIiIiZmZnMzMzMzMy7u7u7u7vMzMzd3d3d3d3d3d27u7u7u7vMzMyqqqqIiIiZmZmIiIh3d3dVVVV3d3eqqqrMzMy7u7u7u7uqqqq7u7u7u7uIiIh3d3eZmZmZmZmZmZmZmZmZmZl3d3dmZmaIiIiZmZmqqqqZmZmZmZm7u7vd3d27u7u7u7uqqqq7u7u7u7uqqqqZmZmIiIiIiIiIiIiIiIh3d3eZmZmIiIiZmZmZmZmqqqqZmZmZmZm7u7vMzMzMzMy7u7uZmZmZmZmqqqqqqqqqqqqqqqqZmZmIiIiZmZm7u7uqqqqqqqq7u7uqqqpmZmZmZmaZmZnMzMzMzMzMzMzMzMy7u7uqqqqIiIiIiIiIiIiZmZmZmZmIiIiZmZmZmZmZmZlmZmaZmZmqqqqZmZmqqqqZmZmIiIh3d3dmZmZmZmZVVVV3d3d3d3dmZmZmZmZ3d3eIiIiZmZl3d3eIiIiZmZmqqqqqqqqqqqqZmZmIiIiZmZmZmZl3d3dmZmaIiIiIiIh3d3eIiIh3d3eIiIiIiIiIiIiqqqqqqqq7u7u7u7u7u7uqqqqqqqqIiIhmZmZ3d3eIiIh3d3eIiIiIiIiIiIiIiIh3d3d3d3eZmZmqqqqZmZm7u7u7u7uqqqq7u7vMzMyZmZmIiIiIiIiZmZmIiIiZmZmZmZmZmZmZmZl3d3dmZmZmZmZmZmZ3d3eZmZmqqqqIiIh3d3dVVVVmZmZmZmZmZmZ3d3eIiIiZmZmZmZmZmZmZmZmZmZmqqqq7u7uIiIhmZmZ3d3eIiIh3d3eIiIh3d3d3d3dVVVVVVVVERERVVVVERERERERVVVVVVVVVVVVmZmZmZmZ3d3d3d3eqqqq7u7uqqqp3d3d3d3d3d3eIiIiIiIh3d3dmZmZVVVVmZmZmZmZ3d3eIiIh3d3d3d3eIiIhVVVVmZmaIiIiZmZmqqqqZmZmIiIiZmZmIiIiIiIh3d3d3d3eZmZmIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3dmZmZVVVV3d3eIiIiqqqqZmZmZmZmIiIh3d3d3d3d3d3dmZmZmZmZ3d3dmZmZVVVVmZmZVVVVVVVVVVVVVVVVERERERERERERVVVV3d3eIiIiZmZl3d3d3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZmZmZVVVVmZmZVVVVEREQzMzMzMzNmZmaIiIiqqqqIiIh3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmaZmZmZmZlVVVVmZmZVVVVERERERERVVVVmZmZVVVVmZmZmZmZmZmZVVVVmZmZmZmZVVVVmZmZmZmZmZmZVVVVmZmZVVVVVVVVVVVVmZmZVVVVVVVVERERERERVVVVmZmZmZmZVVVVmZmZVVVVERERVVVVERERERERERERERERERERERERERERERERVVVVVVVVVVVVEREQzMzMzMzNERERVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERERERVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVVVVVmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3dmZmZVVVVVVVVEREQzMzMzMzMzMzMiIiIiIiJEREREREQiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNVVVVmZmZ3d3dVVVVERERVVVVVVVVERERERERERERERERERERERERERERVVVVVVVVmZmZVVVVVVVVVVVVVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVEREREREQzMzNEREREREREREQzMzMzMzMzMzMzMzNEREQzMzMzMzMiIiIzMzMzMzNERERERERVVVVVVVVVVVVVVVVVVVUzMzMzMzMzMzMzMzNERERVVVVmZmZVVVWIiIi7u7vMzMyIiIhmZmZVVVVVVVV3d3eqqqp3d3czMzNEREQzMzMzMzMzMzMzMzNEREQzMzNEREREREQzMzMzMzMzMzNERERERER3d3eZmZmZmZmZmZl3d3czMzMzMzMzMzMiIiIREREiIiIiIiIzMzMzMzMzMzNEREQzMzMzMzMzMzNERERERERVVVVERERVVVVVVVVERERVVVVVVVVERERVVVVERERVVVVVVVVmZmZVVVVVVVVEREREREREREREREQzMzMzMzMzMzMzMzNERERERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZERERERERERERVVVVVVVVERERERERVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVV3d3d3d3dmZmZVVVVmZmZVVVVVVVVmZmZmZmZVVVVERERVVVVmZmZ3d3dmZmZ3d3d3d3dmZmaZmZm7u7vMzMyqqqpVVVVVVVWZmZl3d3dVVVVVVVVERERmZmZVVVUzMzNEREREREREREREREQzMzNERERERERERERERERVVVVVVVVVVVVmZmZVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVV3d3eIiIiqqqqqqqq7u7vMzMy7u7uZmZlmZmZVVVVVVVVmZmZmZmZVVVUzMzMiIiIzMzMzMzNERERERERVVVVVVVVmZmZVVVVERERERERERERERERERERERERVVVVERERVVVVERERVVVVVVVVVVVVmZmZmZmZERERVVVVVVVVVVVVmZmZmZmZVVVVVVVVmZmZmZmZ3d3d3d3d3d3dmZmZVVVVVVVVVVVVmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZVVVVVVVVERERVVVVVVVV3d3d3d3dmZmZVVVVmZmZ3d3d3d3eIiIiIiIiIiIh3d3d3d3eqqqq7u7vMzMzd3d3d3d3u7u7u7u7MzMyIiIhmZmaqqqqqqqpmZmaIiIiIiIhVVVVERERERERERERVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVEREREREREREREREREREQzMzMzMzMzMzNEREQzMzNERERERERVVVVmZmZVVVUzMzMzMzMzMzNERERVVVV3d3eZmZnMzMzu7u7MzMzMzMzMzMzd3d3u7u7///////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u7u7u7u7u7u7u3d3d3d3dzMzMzMzMzMzMzMzMu7u7zMzMzMzMu7u7zMzMu7u7u7u7zMzMzMzMzMzMu7u7zMzMu7u7u7u7zMzMu7u7u7u7zMzMu7u7zMzMu7u7zMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqmZmZiIiIiIiId3d3d3d3VVVVZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVREREVVVVVVVVREREREREREREREREREREREREREREREREREREREREREREREREMzMzREREREREREREMzMzREREMzMzREREMzMzMzMzMzMzREREMzMzREREREREREREREREMzMzREREMzMzMzMzMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREREREMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREVVVVVVVVREREVVVVREREVVVVZmZmd3d3d3d3ZmZmVVVVVVVVZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmd3d3iIiIiIiIiIiId3d3d3d3d3d3d3d3iIiId3d3ZmZmVVVVZmZmZmZmd3d3d3d3ZmZmREREVVVVVVVVVVVVd3d3u7u7qqqqiIiIiIiImZmZu7u7u7u7u7u7mZmZmZmZd3d3d3d3mZmZzMzM3d3dzMzMu7u73d3d3d3d7u7uzMzMu7u7u7u7u7u7mZmZd3d3iIiIiIiIiIiId3d3d3d3mZmZzMzMzMzMu7u7mZmZmZmZqqqqmZmZiIiImZmZmZmZiIiIiIiIiIiIZmZmd3d3iIiIqqqqqqqqqqqqu7u7u7u7zMzMzMzMu7u7u7u7zMzMu7u7qqqqqqqqmZmZmZmZd3d3iIiIiIiIqqqqqqqqqqqqu7u7u7u7qqqqmZmZiIiIqqqqzMzMu7u7qqqqmZmZmZmZqqqqu7u7qqqqmZmZmZmZqqqqu7u7qqqqqqqqqqqqqqqqmZmZiIiId3d3mZmZu7u7zMzMzMzMu7u7qqqqmZmZmZmZiIiImZmZqqqqiIiIiIiImZmZd3d3ZmZmd3d3qqqqqqqqqqqqqqqqiIiIiIiId3d3ZmZmVVVVZmZmmZmZmZmZiIiIiIiId3d3mZmZd3d3iIiIqqqqqqqqqqqqqqqqmZmZiIiImZmZmZmZd3d3d3d3mZmZmZmZiIiId3d3iIiIiIiId3d3iIiImZmZqqqqqqqqqqqqu7u7qqqqmZmZiIiId3d3d3d3iIiIiIiId3d3iIiIiIiIiIiId3d3d3d3iIiImZmZiIiId3d3iIiImZmZu7u7u7u7qqqqmZmZmZmZmZmZmZmZiIiIiIiIqqqqmZmZd3d3ZmZmZmZmd3d3d3d3iIiIiIiImZmZmZmZd3d3ZmZmd3d3ZmZmd3d3mZmZmZmZmZmZmZmZmZmZmZmZmZmZqqqqd3d3ZmZmiIiIiIiId3d3iIiIiIiIZmZmZmZmZmZmREREVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3mZmZzMzMqqqqmZmZiIiId3d3d3d3d3d3ZmZmZmZmZmZmd3d3d3d3ZmZmd3d3d3d3iIiId3d3ZmZmZmZmiIiImZmZiIiIiIiIiIiImZmZmZmZd3d3ZmZmd3d3iIiIiIiIiIiIiIiIiIiId3d3iIiId3d3iIiIZmZmZmZmiIiIqqqqqqqqiIiIiIiIiIiId3d3d3d3d3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVZmZmVVVVVVVVREREREREREREVVVViIiImZmZmZmZiIiId3d3ZmZmZmZmd3d3ZmZmVVVVVVVVVVVVREREVVVVZmZmZmZmZmZmZmZmREREREREREREVVVVd3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3ZmZmZmZmd3d3mZmZiIiIZmZmZmZmVVVVREREMzMzVVVVZmZmd3d3ZmZmZmZmZmZmVVVVZmZmVVVVZmZmZmZmVVVVZmZmVVVVZmZmVVVVVVVVVVVVZmZmZmZmREREREREREREVVVVZmZmZmZmZmZmZmZmVVVVVVVVREREREREVVVVREREREREREREVVVVREREREREREREVVVVREREREREMzMzREREREREVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREREREREREREREVVVVVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmVVVVZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVREREMzMzREREMzMzIiIiIiIiREREREREMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVVVVVREREVVVVZmZmVVVVREREREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVREREVVVVVVVVREREREREREREREREREREZmZmVVVVREREVVVVZmZmZmZmVVVVREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREVVVVREREVVVVVVVVVVVVREREMzMzMzMzIiIiMzMzVVVVVVVVVVVVVVVVd3d3u7u7u7u7iIiIVVVVVVVVREREZmZmiIiIVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzMzMzMzMzREREREREiIiImZmZmZmZmZmZd3d3VVVVREREMzMzMzMzMzMzIiIiIiIiMzMzMzMzREREREREREREREREMzMzMzMzREREREREVVVVREREREREVVVVREREVVVVREREVVVVVVVVVVVVZmZmVVVVZmZmREREREREMzMzMzMzREREMzMzMzMzMzMzREREREREREREREREREREREREZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREVVVVREREREREVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmd3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVd3d3iIiId3d3d3d3iIiIZmZmd3d3qqqqzMzMqqqqREREVVVVmZmZZmZmVVVVREREVVVVZmZmVVVVREREREREREREREREMzMzREREREREREREVVVVREREVVVVZmZmVVVVVVVVZmZmVVVVREREVVVVVVVVVVVVREREVVVVZmZmVVVVd3d3mZmZmZmZqqqqu7u7u7u7qqqqiIiIZmZmZmZmZmZmZmZmVVVVREREMzMzMzMzMzMzREREREREREREVVVVZmZmZmZmVVVVREREREREREREREREREREVVVVVVVVVVVVREREVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVZmZmd3d3d3d3d3d3d3d3iIiIqqqqqqqqmZmZiIiImZmZiIiImZmZu7u73d3d7u7u7u7u3d3dqqqqiIiImZmZd3d3VVVVZmZmiIiIZmZmZmZmVVVVVVVVREREVVVVVVVVZmZmZmZmVVVVVVVVVVVVZmZmd3d3ZmZmREREREREREREREREMzMzMzMzREREMzMzMzMzMzMzREREVVVVVVVVVVVVMzMzMzMzMzMzREREMzMzREREVVVViIiIqqqq3d3d3d3dzMzMu7u73d3d7u7u////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7szMzLu7u6qqqpmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiJmZmYiIiJmZmYiIiHd3d4iIiIiIiIiIiIiIiJmZmZmZmaqqqqqqqqqqqqqqqru7u6qqqru7u7u7u6qqqqqqqqqqqqqqqpmZmaqqqpmZmYiIiIiIiHd3d2ZmZlVVVVVVVURERERERERERERERERERERERERERERERDMzM0RERERERDMzMzMzM0RERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIhERESIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIjMzMyIiIiIiIjMzMyIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzM0RERERERERERFVVVURERERERERERFVVVWZmZmZmZmZmZmZmZlVVVWZmZnd3d4iIiGZmZmZmZnd3d5mZmXd3d1VVVVVVVWZmZoiIiIiIiIiIiHd3d3d3d4iIiJmZmYiIiIiIiHd3d2ZmZmZmZlVVVVVVVWZmZmZmZmZmZlVVVVVVVURERFVVVYiIiKqqqqqqqnd3d2ZmZnd3d6qqqru7u5mZmYiIiJmZmZmZmYiIiJmZmczMzN3d3d3d3d3d3d3d3e7u7t3d3czMzLu7u7u7u6qqqpmZmXd3d3d3d4iIiIiIiIiIiIiIiJmZmczMzN3d3aqqqqqqqpmZmYiIiIiIiJmZmZmZmZmZmZmZmXd3d2ZmZnd3d4iIiKqqqru7u6qqqqqqqru7u6qqqru7u8zMzMzMzLu7u8zMzLu7u7u7u6qqqpmZmZmZmYiIiHd3d5mZmbu7u8zMzLu7u7u7u6qqqqqqqoiIiHd3d5mZmbu7u7u7u5mZmaqqqpmZmaqqqpmZmXd3d4iIiKqqqru7u6qqqpmZmaqqqqqqqpmZmZmZmbu7u4iIiHd3d6qqqru7u7u7u7u7u6qqqqqqqpmZmYiIiJmZmaqqqoiIiHd3d4iIiIiIiGZmZnd3d5mZmaqqqqqqqqqqqqqqqoiIiIiIiGZmZmZmZoiIiJmZmZmZmZmZmYiIiIiIiIiIiIiIiJmZmaqqqpmZmZmZmZmZmaqqqpmZmZmZmZmZmYiIiJmZmZmZmZmZmZmZmYiIiIiIiIiIiIiIiIiIiJmZmaqqqpmZmYiIiJmZmaqqqoiIiJmZmZmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d4iIiIiIiGZmZnd3d6qqqszMzLu7u5mZmbu7u6qqqpmZmaqqqpmZmZmZmaqqqpmZmXd3d3d3d3d3d4iIiIiIiHd3d3d3d4iIiJmZmXd3d3d3d2ZmZnd3d3d3d5mZmZmZmZmZmZmZmZmZmaqqqpmZmYiIiIiIiJmZmaqqqmZmZmZmZpmZmYiIiGZmZmZmZlVVVURERFVVVURERFVVVURERFVVVVVVVWZmZmZmZmZmZnd3d6qqqru7u7u7u5mZmYiIiHd3d2ZmZmZmZmZmZnd3d3d3d4iIiHd3d3d3d3d3d2ZmZnd3d4iIiGZmZmZmZoiIiJmZmYiIiIiIiHd3d4iIiIiIiIiIiHd3d3d3d4iIiIiIiJmZmZmZmYiIiIiIiIiIiIiIiIiIiGZmZmZmZpmZmbu7u6qqqpmZmYiIiIiIiHd3d3d3d3d3d2ZmZlVVVWZmZmZmZlVVVVVVVWZmZmZmZlVVVVVVVURERDMzM0RERFVVVYiIiJmZmaqqqpmZmYiIiGZmZmZmZmZmZlVVVWZmZlVVVVVVVURERFVVVVVVVWZmZmZmZlVVVVVVVVVVVURERFVVVXd3d4iIiHd3d4iIiIiIiHd3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZnd3d4iIiHd3d1VVVVVVVVVVVURERDMzM0RERGZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZlVVVWZmZmZmZlVVVVVVVURERERERERERGZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVURERERERERERERERERERERERERERDMzM0RERERERERERDMzMzMzM0RERGZmZmZmZlVVVWZmZmZmZmZmZlVVVWZmZlVVVURERERERERERERERFVVVURERERERERERERERERERERERERERFVVVVVVVURERGZmZmZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZlVVVVVVVURERERERDMzMzMzMzMzMzMzMyIiIkRERERERDMzMyIiIiIiIjMzMyIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVURERDMzM0RERERERERERFVVVVVVVVVVVVVVVURERFVVVURERERERERERERERERERERERERERERERERERERERERERERERERERERERFVVVWZmZkRERFVVVVVVVWZmZlVVVVVVVURERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzM0RERFVVVVVVVVVVVVVVVURERDMzMzMzMzMzMyIiIjMzM0RERFVVVWZmZmZmZoiIiMzMzKqqqmZmZlVVVVVVVURERGZmZnd3d0RERERERDMzMzMzMyIiIjMzMzMzMzMzM0RERFVVVURERDMzMyIiIjMzMzMzM0RERHd3d6qqqqqqqpmZmYiIiGZmZlVVVURERERERERERDMzMyIiIjMzMzMzMzMzM1VVVURERERERDMzM0RERERERERERERERFVVVURERERERFVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVURERDMzM0RERDMzM0RERDMzM0RERERERERERERERERERERERFVVVVVVVWZmZlVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERFVVVURERFVVVWZmZkRERFVVVVVVVVVVVVVVVVVVVURERFVVVVVVVWZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmaqqqoiIiIiIiIiIiGZmZnd3d5mZmczMzIiIiDMzM1VVVZmZmWZmZlVVVVVVVVVVVWZmZkRERERERERERDMzM0RERERERDMzM0RERERERFVVVVVVVVVVVVVVVVVVVURERFVVVURERERERFVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZoiIiJmZmZmZmbu7u7u7u5mZmaqqqpmZmWZmZmZmZmZmZmZmZmZmZjMzMzMzMzMzM0RERERERERERERERFVVVWZmZlVVVVVVVURERERERERERFVVVVVVVURERERERFVVVURERFVVVVVVVVVVVVVVVXd3d4iIiHd3d1VVVWZmZmZmZlVVVWZmZlVVVVVVVWZmZlVVVWZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVURERFVVVWZmZmZmZmZmZlVVVXd3d3d3d4iIiJmZmXd3d5mZmaqqqqqqqoiIiHd3d5mZmZmZmZmZmZmZmczMzN3d3e7u7t3d3czMzJmZmWZmZmZmZmZmZoiIiJmZmXd3d1VVVVVVVVVVVURERERERERERGZmZlVVVVVVVURERFVVVWZmZoiIiIiIiGZmZlVVVURERERERDMzMzMzMzMzMzMzM0RERDMzM0RERFVVVVVVVTMzMzMzMyIiIjMzMzMzMzMzM0RERFVVVXd3d5mZmbu7u93d3bu7u8zMzMzMzO7u7u7u7v///////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7d3d3d3d3MzMy7u7u7u7vMzMzMzMy7u7u7u7u7u7vMzMy7u7u7u7uqqqqqqqqZmZmqqqqZmZmIiIiZmZmIiIiZmZmZmZmqqqq7u7u7u7vMzMzMzMzMzMzd3d3MzMzd3d3MzMzd3d3d3d3d3d3MzMzMzMzMzMzMzMzMzMy7u7uqqqqqqqqZmZmZmZmIiIiIiIiIiIh3d3eIiIh3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVmZmZmZmZVVVVEREREREREREREREREREREREQzMzNEREREREREREREREREREQzMzMzMzMzMzNEREREREREREQzMzMzMzMzMzNEREREREQzMzNEREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMiIiIiIiIiIiIiIiIzMzMzMzNEREREREQzMzMzMzMzMzMzMzNERERERERERERVVVVVVVVERERERERVVVVVVVVmZmZVVVVmZmZVVVVmZmZmZmZVVVVmZmZmZmaIiIiZmZmZmZmIiIh3d3d3d3d3d3d3d3d3d3d3d3eIiIiZmZmZmZmZmZl3d3d3d3dmZmZVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVUzMzNVVVWZmZnMzMyqqqp3d3dERER3d3eIiIiZmZmIiIiIiIiqqqrMzMy7u7uqqqq7u7vd3d3u7u7d3d3d3d3d3d3d3d3d3d3MzMy7u7uZmZmIiIiZmZmZmZmZmZmZmZmZmZmZmZmZmZm7u7u7u7u7u7uqqqqZmZl3d3eZmZmZmZmZmZl3d3d3d3dVVVVmZmZmZmaqqqrMzMy7u7u7u7uqqqq7u7uqqqqqqqq7u7vMzMzMzMy7u7u7u7vMzMyqqqqIiIiIiIiIiIhmZmaIiIi7u7vd3d27u7uqqqqqqqqZmZl3d3dmZmaIiIiqqqq7u7u7u7u7u7uqqqq7u7uqqqp3d3d3d3e7u7uqqqqIiIiIiIiqqqq7u7uqqqqZmZmZmZmZmZlmZmZ3d3eZmZm7u7u7u7uqqqqqqqqZmZmZmZmZmZmqqqqZmZmIiIhmZmaIiIiIiIh3d3eIiIiZmZmZmZmIiIiIiIiZmZmZmZmIiIiIiIiZmZmZmZmIiIiqqqqZmZmIiIiZmZmIiIiIiIiZmZmZmZmZmZmIiIiZmZmZmZmZmZmIiIiZmZmZmZmIiIiZmZmZmZmIiIiIiIiIiIiIiIiIiIiqqqqqqqqIiIiIiIiIiIiIiIiZmZmZmZmqqqqZmZmZmZmZmZmIiIiIiIiIiIiIiIiIiIh3d3eIiIiIiIiIiIhmZmZmZmaZmZnMzMy7u7u7u7u7u7uqqqqqqqqqqqqqqqqqqqq7u7uZmZmIiIh3d3eIiIiIiIiIiIh3d3d3d3eIiIiZmZmIiIh3d3d3d3dmZmaIiIiIiIiZmZmZmZmZmZmZmZmIiIiIiIiZmZmZmZmqqqqZmZl3d3eIiIiqqqp3d3dERERVVVVmZmZVVVVERERVVVVERERERERERERVVVVVVVVVVVVVVVVmZmaZmZnMzMy7u7uZmZl3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3d3d3dmZmaIiIh3d3dmZmZmZmZ3d3eZmZmIiIiIiIh3d3eIiIiIiIiIiIiIiIh3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIhmZmZVVVWIiIiZmZmqqqqZmZmIiIh3d3d3d3dmZmZmZmZmZmZVVVVmZmZmZmZmZmZVVVVVVVVmZmZmZmZEREREREQzMzNERERERER3d3eIiIiqqqqZmZmZmZmIiIhmZmZmZmZVVVVVVVVVVVVERERERERERERVVVVmZmZVVVVmZmZmZmZVVVVERERERER3d3eIiIiIiIiIiIh3d3dmZmZmZmZmZmZ3d3dmZmZmZmZVVVVVVVVVVVV3d3d3d3dmZmZmZmZmZmZVVVVERERVVVVVVVVmZmZmZmZmZmZ3d3dVVVVmZmZmZmZVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVERERVVVVEREREREREREQzMzNVVVVVVVVmZmZmZmZmZmZVVVVVVVVEREREREQzMzNEREQzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzNEREREREREREQzMzMzMzNmZmZVVVVmZmZmZmZ3d3dmZmZVVVVmZmZERERVVVVERERERERVVVVEREQzMzNEREQzMzNERERVVVVERERERERVVVVERERERERVVVVmZmZERERVVVVVVVVmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVEREREREQzMzMzMzMiIiIzMzMiIiIiIiJERERVVVUzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIzMzMzMzMzMzNEREQzMzMzMzMiIiJERERVVVVmZmZmZmZmZmZVVVVERERVVVVERERERERVVVVVVVVEREREREREREREREREREREREQzMzNERERERERERERVVVVVVVVERERVVVVERERVVVVVVVVVVVVEREREREREREREREREREQzMzMzMzNEREREREQzMzMzMzMzMzMzMzNEREQzMzNERERERERVVVVVVVVVVVVEREREREREREQzMzMzMzMzMzMzMzNVVVVmZmaIiIiqqqq7u7uIiIhERERERERERERmZmaIiIhmZmZEREQzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERVVVVEREQzMzMzMzMzMzMzMzNERESZmZmqqqqZmZmIiIiIiIhmZmZVVVVEREREREQiIiIREREiIiIzMzNEREREREREREREREREREQzMzNERERERERERERERERVVVVERERVVVVERERERERERERVVVVVVVVVVVVVVVVERERERERERERERERERERERERERERERERERERVVVVVVVVmZmZERERERERERERERERERERERERVVVVVVVVVVVVERERVVVVERERERERERERERERVVVVVVVVERERVVVVVVVVERERERERERERVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVERERVVVVVVVV3d3eZmZl3d3dmZmZmZmZVVVVmZmaZmZnMzMx3d3czMzNVVVWZmZl3d3dmZmZmZmZVVVVmZmZVVVVEREREREREREQzMzNERERERERERERERERERERERERERERVVVVVVVVVVVVERERERERERERVVVVmZmZ3d3eIiIhmZmZmZmZVVVVERERVVVWIiIiZmZm7u7uqqqqZmZmIiIiZmZmIiIh3d3dmZmZ3d3dmZmZmZmZVVVVERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVV3d3d3d3d3d3dmZmZmZmZmZmZVVVVVVVVERERVVVVVVVVERERVVVVERERERERmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZVVVVERERERERERERERERVVVVmZmZmZmZVVVVmZmZmZmZ3d3d3d3d3d3d3d3eqqqqqqqqIiIhmZmaIiIiIiIiqqqq7u7u7u7u7u7u7u7vMzMzMzMyZmZl3d3dVVVV3d3eIiIiIiIhmZmZ3d3d3d3d3d3dmZmZERERERERERERERERVVVVERERVVVVmZmZ3d3eIiIh3d3dmZmZVVVVEREREREQzMzMzMzNEREQzMzNERERVVVVEREREREQzMzMiIiIzMzMzMzNEREQzMzNERERVVVVVVVVmZmaZmZnMzMzMzMy7u7u7u7vd3d3///////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////3d3d3d3d3d3d7u7u3d3d3d3d3d3d7u7u7u7u7u7u3d3d3d3d3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzMzMzM3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3dzMzMzMzMu7u7u7u7qqqqqqqqqqqqmZmZmZmZmZmZmZmZiIiImZmZmZmZmZmZmZmZqqqqmZmZqqqqqqqqqqqqmZmZmZmZiIiIiIiImZmZiIiId3d3iIiId3d3ZmZmd3d3d3d3ZmZmZmZmd3d3ZmZmZmZmd3d3ZmZmVVVVVVVVVVVVVVVVVVVVREREREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVREREVVVVREREREREREREREREMzMzREREREREMzMzREREREREMzMzMzMzMzMzMzMzREREMzMzREREREREREREREREREREMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiMzMzMzMzMzMzREREREREREREMzMzMzMzREREREREVVVVVVVVVVVVZmZmd3d3VVVVd3d3d3d3ZmZmZmZmZmZmd3d3d3d3ZmZmVVVVMzMzVVVViIiImZmZqqqqmZmZmZmZmZmZd3d3ZmZmZmZmZmZmiIiImZmZmZmZmZmZiIiId3d3ZmZmZmZmZmZmVVVVd3d3ZmZmVVVVVVVVVVVVREREREREd3d3u7u7zMzMqqqqd3d3ZmZmd3d3iIiIiIiImZmZqqqqu7u7zMzMu7u7qqqqu7u77u7u3d3d3d3d3d3dzMzM3d3d7u7u3d3du7u7mZmZiIiImZmZmZmZqqqqmZmZqqqqmZmZqqqqqqqqqqqqu7u7mZmZiIiIiIiImZmZqqqqiIiIVVVVVVVVVVVVVVVVd3d3qqqqu7u7u7u7u7u7qqqqqqqqmZmZqqqqu7u7zMzMu7u7qqqqqqqqqqqqmZmZiIiIiIiIiIiIiIiImZmZzMzMzMzMqqqqqqqqqqqqqqqqiIiIiIiImZmZqqqqu7u7zMzMu7u7zMzMu7u7iIiId3d3qqqqu7u7mZmZiIiImZmZu7u7u7u7qqqqmZmZmZmZmZmZd3d3ZmZmiIiImZmZu7u7qqqqqqqqqqqqqqqqu7u7qqqqqqqqmZmZd3d3ZmZmiIiIiIiIiIiImZmZmZmZZmZmd3d3iIiImZmZmZmZqqqqmZmZd3d3iIiImZmZmZmZqqqqqqqqiIiIiIiIiIiImZmZmZmZZmZmd3d3mZmZiIiIiIiIqqqqu7u7mZmZiIiIiIiIiIiImZmZmZmZmZmZmZmZmZmZqqqqiIiIiIiId3d3iIiImZmZqqqqmZmZqqqqqqqqmZmZiIiIiIiIiIiImZmZiIiIiIiId3d3iIiId3d3ZmZmd3d3qqqqzMzMzMzMqqqqu7u7qqqqiIiIiIiImZmZqqqqu7u7mZmZmZmZmZmZiIiIiIiIiIiIiIiIZmZmiIiImZmZmZmZd3d3ZmZmd3d3d3d3iIiImZmZiIiIiIiIiIiIiIiId3d3iIiImZmZqqqqmZmZiIiIiIiIu7u7ZmZmVVVVVVVVREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmmZmZzMzMu7u7mZmZiIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3iIiId3d3ZmZmVVVVd3d3mZmZiIiIiIiIiIiImZmZiIiIiIiIiIiIiIiId3d3iIiId3d3d3d3iIiIiIiIiIiIiIiIiIiIVVVVVVVVd3d3mZmZqqqqmZmZd3d3ZmZmZmZmd3d3ZmZmVVVVVVVVREREZmZmZmZmZmZmZmZmZmZmZmZmVVVVREREMzMzREREMzMzZmZmiIiImZmZiIiIiIiId3d3d3d3VVVVVVVVVVVVREREREREREREVVVVZmZmZmZmZmZmVVVVZmZmVVVVMzMzVVVVZmZmiIiId3d3d3d3iIiIVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVZmZmd3d3d3d3ZmZmVVVVZmZmVVVVVVVVREREVVVVZmZmZmZmZmZmVVVVZmZmREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREVVVVVVVVREREMzMzMzMzVVVVVVVVVVVVZmZmVVVVVVVVMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzREREREREREREREREMzMzMzMzREREVVVVVVVVZmZmd3d3VVVVREREREREMzMzREREVVVVREREREREREREMzMzREREMzMzMzMzREREREREVVVVVVVVMzMzREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVREREVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVREREMzMzMzMzIiIiIiIiIiIiIiIiMzMzREREVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzREREREREMzMzMzMzREREZmZmVVVVZmZmZmZmVVVVVVVVREREREREVVVVVVVVREREVVVVREREREREREREREREREREREREREREREREREREREREREREREREVVVVREREREREREREREREREREREREREREREREMzMzREREMzMzMzMzMzMzREREMzMzMzMzREREREREMzMzMzMzMzMzREREVVVVREREREREREREREREMzMzREREMzMzREREREREVVVVd3d3mZmZmZmZZmZmREREMzMzVVVVmZmZiIiIVVVVMzMzREREMzMzMzMzMzMzMzMzREREREREREREREREREREREREMzMzIiIiMzMzREREREREZmZmmZmZiIiImZmZiIiIZmZmVVVVREREIiIiIiIiIiIiERERIiIiMzMzMzMzREREREREREREREREREREREREVVVVVVVVREREVVVVREREREREREREVVVVVVVVVVVVVVVVREREREREREREREREREREREREVVVVVVVVVVVVREREREREVVVVZmZmVVVVREREREREREREREREREREVVVVVVVVVVVVVVVVREREREREREREREREREREVVVVVVVVREREREREVVVVVVVVVVVVREREVVVVVVVVVVVVREREZmZmZmZmZmZmZmZmZmZmVVVVVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVZmZmqqqqu7u7ZmZmMzMzVVVViIiIiIiId3d3VVVVVVVVZmZmVVVVREREREREREREREREREREREREVVVVREREMzMzREREREREVVVVVVVVVVVVREREREREVVVVVVVVVVVVZmZmd3d3ZmZmZmZmVVVVREREVVVVZmZmiIiImZmZqqqqmZmZiIiId3d3iIiId3d3d3d3ZmZmd3d3d3d3d3d3d3d3ZmZmVVVVREREREREREREREREREREVVVVZmZmVVVVZmZmZmZmZmZmVVVVVVVVZmZmVVVVZmZmVVVVZmZmZmZmZmZmd3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVZmZmd3d3d3d3ZmZmZmZmZmZmVVVVZmZmZmZmVVVVREREREREMzMzVVVVVVVVZmZmVVVVVVVVZmZmd3d3d3d3d3d3ZmZmZmZmqqqqu7u7mZmZiIiId3d3d3d3mZmZzMzMu7u7qqqqiIiIqqqqmZmZqqqqmZmZd3d3d3d3ZmZmZmZmd3d3mZmZiIiIZmZmZmZmVVVVREREMzMzREREREREREREREREVVVVZmZmVVVVZmZmVVVVREREREREREREREREMzMzMzMzREREREREREREREREMzMzIiIiMzMzMzMzMzMzMzMzREREREREVVVVVVVVVVVVd3d3qqqqzMzMzMzMqqqqzMzM7u7u////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7t3d3d3d3d3d3e7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3d3d3d3d3e7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3czMzMzMzLu7u6qqqpmZmZmZmYiIiJmZmZmZmYiIiJmZmYiIiIiIiIiIiJmZmYiIiJmZmZmZmaqqqqqqqqqqqqqqqqqqqqqqqpmZmZmZmZmZmZmZmZmZmZmZmZmZmYiIiJmZmZmZmYiIiJmZmYiIiIiIiJmZmZmZmYiIiIiIiIiIiHd3d3d3d2ZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVWZmZlVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVURERERERERERERERERERERERFVVVURERERERERERERERERERERERFVVVURERERERFVVVURERERERERERERERDMzMzMzM0RERERERERERERERDMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERFVVVVVVVVVVVWZmZnd3d5mZmYiIiHd3d3d3d4iIiHd3d3d3d3d3d4iIiHd3d1VVVURERERERGZmZoiIiJmZmZmZmZmZmZmZmZmZmYiIiHd3d2ZmZmZmZpmZmZmZmZmZmZmZmYiIiGZmZmZmZnd3d2ZmZmZmZnd3d2ZmZmZmZlVVVURERDMzM0RERGZmZqqqqszMzKqqqoiIiHd3d2ZmZnd3d4iIiKqqqru7u8zMzLu7u7u7u5mZmZmZmczMzN3d3czMzMzMzN3d3d3d3d3d3d3d3czMzJmZmYiIiIiIiKqqqpmZmZmZmZmZmZmZmaqqqpmZmaqqqpmZmZmZmXd3d4iIiKqqqpmZmVVVVVVVVURERFVVVVVVVZmZmaqqqqqqqqqqqqqqqru7u6qqqpmZmaqqqru7u7u7u7u7u6qqqqqqqpmZmZmZmYiIiJmZmaqqqru7u8zMzMzMzLu7u6qqqru7u7u7u6qqqru7u6qqqpmZmZmZmaqqqqqqqqqqqru7u7u7u4iIiIiIiLu7u7u7u5mZmYiIiJmZmbu7u8zMzKqqqqqqqpmZmaqqqpmZmXd3d3d3d4iIiIiIiJmZmZmZmaqqqru7u7u7u6qqqpmZmYiIiIiIiHd3d3d3d3d3d4iIiJmZmXd3d3d3d3d3d4iIiHd3d5mZmaqqqqqqqoiIiJmZmYiIiJmZmZmZmZmZmYiIiIiIiIiIiIiIiIiIiGZmZlVVVVVVVXd3d6qqqszMzKqqqqqqqoiIiJmZmaqqqqqqqqqqqpmZmZmZmZmZmZmZmYiIiIiIiHd3d5mZmaqqqqqqqqqqqqqqqru7u6qqqpmZmZmZmYiIiHd3d4iIiIiIiGZmZmZmZmZmZnd3d3d3d5mZmczMzMzMzKqqqqqqqqqqqpmZmYiIiIiIiKqqqru7u6qqqqqqqqqqqqqqqpmZmZmZmYiIiHd3d5mZmaqqqqqqqoiIiGZmZmZmZnd3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiJmZmYiIiHd3d3d3d7u7u4iIiFVVVURERDMzMzMzMzMzM1VVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVXd3d5mZmczMzLu7u6qqqoiIiHd3d3d3d3d3d3d3d4iIiHd3d3d3d4iIiHd3d3d3d3d3d5mZmXd3d1VVVVVVVXd3d5mZmYiIiJmZmYiIiIiIiJmZmYiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiJmZmYiIiHd3d2ZmZlVVVXd3d4iIiJmZmZmZmXd3d3d3d3d3d3d3d2ZmZlVVVURERERERFVVVXd3d2ZmZmZmZmZmZlVVVURERERERDMzMzMzMzMzM1VVVZmZmaqqqoiIiIiIiHd3d2ZmZmZmZlVVVURERERERERERFVVVURERGZmZmZmZmZmZmZmZkRERERERDMzM0RERGZmZoiIiIiIiIiIiHd3d2ZmZlVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVWZmZmZmZlVVVVVVVVVVVURERFVVVURERFVVVXd3d2ZmZlVVVVVVVVVVVVVVVURERERERERERFVVVVVVVWZmZlVVVURERFVVVURERFVVVURERERERERERERERERERFVVVWZmZlVVVVVVVVVVVURERDMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERERERFVVVURERDMzMzMzM1VVVVVVVVVVVWZmZlVVVVVVVURERDMzMzMzM0RERERERERERDMzMzMzM0RERDMzM0RERERERERERFVVVVVVVURERDMzMzMzM1VVVWZmZlVVVVVVVWZmZmZmZlVVVURERERERERERERERFVVVURERERERERERERERERERERERFVVVVVVVURERDMzMzMzMzMzMzMzMyIiIiIiIjMzM0RERERERERERERERDMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMyIiIiIiIhERESIiIiIiIiIiIiIiIjMzM0RERERERERERERERERERERERFVVVVVVVVVVVWZmZlVVVVVVVURERFVVVVVVVVVVVURERERERERERERERDMzM0RERDMzM0RERERERERERERERFVVVURERERERERERERERFVVVVVVVURERFVVVURERDMzM0RERERERDMzM0RERDMzMzMzMzMzM0RERERERERERDMzMzMzMzMzM0RERDMzM0RERERERERERDMzMzMzM0RERDMzM0RERERERERERERERFVVVYiIiIiIiFVVVURERERERHd3d5mZmWZmZkRERERERDMzMzMzM1VVVURERDMzM0RERERERERERFVVVVVVVVVVVTMzMzMzMzMzM0RERERERGZmZnd3d5mZmaqqqoiIiHd3d2ZmZkRERCIiIiIiIiIiIhERESIiIjMzMzMzMzMzM0RERFVVVURERERERFVVVVVVVURERFVVVVVVVVVVVVVVVURERGZmZmZmZmZmZlVVVVVVVVVVVURERERERERERFVVVVVVVURERERERERERFVVVVVVVVVVVURERERERERERERERERERERERERERFVVVVVVVVVVVURERERERERERERERFVVVVVVVVVVVURERFVVVURERFVVVVVVVURERFVVVVVVVVVVVVVVVWZmZnd3d2ZmZmZmZmZmZlVVVURERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZkRERHd3d6qqqpmZmURERDMzM1VVVaqqqpmZmXd3d2ZmZlVVVWZmZlVVVVVVVURERFVVVURERERERERERERERERERERERERERFVVVVVVVURERFVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZlVVVVVVVVVVVURERERERFVVVXd3d5mZmZmZmaqqqpmZmZmZmXd3d3d3d3d3d4iIiHd3d3d3d3d3d4iIiIiIiGZmZmZmZlVVVURERERERERERERERFVVVVVVVVVVVWZmZlVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZlVVVWZmZlVVVVVVVURERFVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZlVVVVVVVURERERERDMzM1VVVWZmZlVVVURERFVVVWZmZmZmZqqqqoiIiGZmZmZmZpmZmbu7u7u7u4iIiJmZmXd3d3d3d4iIiKqqqpmZmZmZmaqqqqqqqqqqqru7u3d3d2ZmZmZmZmZmZmZmZoiIiIiIiGZmZlVVVURERERERDMzM0RERERERERERERERERERERERERERFVVVVVVVURERERERERERERERERERDMzM0RERERERERERERERCIiIjMzMyIiIjMzMzMzM0RERERERERERFVVVVVVVVVVVXd3d4iIiLu7u8zMzLu7u8zMzO7u7v///////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////u7u7d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3MzMy7u7vMzMzMzMzMzMzMzMy7u7vMzMzd3d3MzMzd3d3d3d3d3d3u7u7d3d3u7u7d3d3u7u7u7u7u7u7d3d3u7u7d3d3u7u7d3d3d3d3d3d3d3d3MzMzMzMy7u7uqqqqqqqqqqqqZmZmZmZmZmZmZmZmZmZmIiIiIiIiIiIiIiIiZmZmIiIiIiIiqqqqqqqqZmZmIiIiZmZmZmZmZmZmIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIiIiIiIiIiZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIiIiIh3d3d3d3eIiIh3d3eIiIh3d3d3d3d3d3d3d3eIiIh3d3d3d3d3d3dmZmZmZmZmZmZVVVVmZmZVVVVVVVVVVVVmZmZVVVVVVVVVVVVERERVVVVVVVVERERERERVVVVEREREREREREQzMzNEREREREQzMzMzMzNEREQzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREREREQzMzMzMzNEREQzMzNERERVVVVVVVVmZmZ3d3eZmZl3d3dmZmZ3d3eIiIiZmZmIiIiZmZmIiIhVVVVVVVVmZmZmZmZmZmZ3d3d3d3dmZmZ3d3eIiIiZmZmIiIhmZmZVVVVmZmaIiIiZmZmIiIiZmZmIiIhmZmZmZmZ3d3d3d3dmZmZVVVVmZmZmZmZEREREREQzMzNERERmZmaqqqrMzMyqqqqIiIh3d3dmZmZ3d3eqqqrMzMzMzMy7u7u7u7u7u7uZmZmZmZm7u7vMzMzMzMzMzMzd3d3d3d3MzMzMzMy7u7uqqqp3d3eZmZmqqqqZmZmIiIiIiIiZmZm7u7uqqqqZmZmIiIiIiIiIiIiZmZm7u7t3d3dVVVVERERERERERER3d3eqqqqqqqqqqqqqqqq7u7u7u7uqqqqqqqq7u7uqqqqqqqq7u7u7u7uqqqqZmZmZmZmIiIiqqqrMzMzMzMzd3d3MzMyqqqq7u7vMzMy7u7u7u7u7u7uqqqqZmZmZmZmqqqqqqqqqqqqZmZmZmZmIiIiqqqrMzMy7u7uIiIiIiIiZmZmqqqq7u7uqqqqqqqqqqqq7u7uqqqqZmZl3d3d3d3eIiIh3d3eZmZm7u7vMzMy7u7uqqqqZmZmIiIiZmZmZmZmIiIhmZmZ3d3eIiIiIiIh3d3dmZmZVVVVVVVWIiIi7u7uqqqqIiIiZmZmqqqqZmZmZmZmZmZmZmZmIiIh3d3d3d3dmZmZ3d3dVVVVERESIiIi7u7vMzMy7u7uqqqqZmZmqqqqqqqqqqqqqqqqZmZmqqqqZmZmZmZmZmZl3d3d3d3eZmZmqqqqqqqqqqqqqqqq7u7uqqqqZmZmZmZmIiIiIiIiZmZmIiIhmZmZmZmZmZmZmZmZmZmaIiIjMzMyqqqqqqqqqqqqqqqqZmZl3d3d3d3eqqqqqqqqqqqq7u7u7u7uqqqqZmZmZmZmZmZmZmZmZmZmqqqqZmZmZmZl3d3d3d3dmZmZ3d3dmZmZ3d3eIiIiIiIiIiIh3d3eIiIiZmZmIiIh3d3dVVVV3d3eZmZlmZmZVVVVEREQzMzMzMzMzMzNERERVVVVVVVVVVVVERERmZmZmZmZVVVV3d3eZmZm7u7u7u7uqqqqIiIiIiIh3d3d3d3d3d3d3d3eIiIh3d3d3d3dmZmZ3d3eIiIh3d3dmZmZVVVVmZmaIiIiZmZmZmZmZmZmIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3dmZmaIiIiIiIiZmZl3d3dmZmZmZmZVVVVmZmZ3d3eZmZmqqqqIiIh3d3d3d3dmZmZVVVVVVVVERERERERmZmZ3d3dmZmZmZmZmZmZVVVVVVVVEREQzMzMzMzMiIiJERESZmZmqqqqZmZl3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVmZmZmZmZVVVVEREQzMzNERERERERVVVV3d3eIiIh3d3eIiIhmZmZERERERERVVVVmZmZmZmZmZmZVVVVmZmZ3d3dVVVVERERERERERERVVVVVVVVERERVVVVmZmZmZmZVVVVVVVVVVVVVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVERERVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNEREREREREREREREREREQzMzNERERERERERERVVVVmZmZVVVVVVVVEREQzMzMzMzNEREQzMzMzMzMzMzMzMzNEREQzMzNERERERERERERVVVVVVVVVVVUzMzMzMzNERERVVVV3d3dmZmZVVVVmZmZVVVVERERERERERERERERVVVVERERERERVVVVEREREREREREQzMzNEREREREREREREREREREQzMzMzMzMzMzMzMzNEREREREQzMzNEREREREQzMzMiIiIzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzNEREQzMzNERERVVVVERERERERERERERERVVVVVVVVVVVVERERERERERERERERERERVVVVEREQzMzNEREREREQzMzNERERERERERERVVVVVVVVERERERERERERERERERERmZmZVVVVERERERERVVVVEREREREREREREREQzMzMzMzNEREQzMzNEREREREQzMzNEREQzMzMzMzNEREREREREREQzMzNEREREREQzMzNERERERERERERVVVVERERERERERERmZmZmZmZVVVVERERERESIiIiIiIhVVVVEREQzMzNERERERERERERVVVVERERERERVVVVVVVVVVVVmZmZVVVVEREQzMzMiIiIzMzNERERmZmaIiIiqqqqqqqqZmZl3d3dVVVVEREQzMzMiIiIREREiIiIREREiIiIzMzNERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVmZmZmZmZERERERERVVVVERERERERERERERERERERERERERERERERVVVVEREREREREREREREREREREREREREREREQzMzNERERVVVVVVVVVVVVERERERERERERERERVVVVVVVVERERVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVmZmZ3d3d3d3dmZmZERERERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVV3d3dmZmZVVVVVVVV3d3e7u7uIiIgzMzMiIiJmZma7u7uqqqp3d3dmZmZVVVVmZmZVVVVVVVVVVVVERERERERERERERERERERERERERERERERERERVVVVERERERERVVVVVVVVmZmZmZmZ3d3d3d3d3d3d3d3dmZmZVVVVERERVVVVVVVVmZmZ3d3eZmZmZmZmZmZmZmZmIiIiIiIiIiIiIiIiIiIh3d3d3d3eIiIh3d3d3d3d3d3dmZmZmZmZVVVVERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVmZmZmZmZ3d3eIiIh3d3dmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZVVVVmZmZmZmZmZmZVVVVERERVVVVERERERERmZmZ3d3dVVVVERERVVVVVVVVmZmaIiIiZmZlmZmZVVVV3d3e7u7u7u7uZmZmIiIh3d3dmZmaIiIiZmZmqqqqZmZmZmZmZmZmqqqqqqqqIiIhVVVVmZmZmZmZmZmZmZmZ3d3eIiIh3d3dVVVVERERERERVVVVEREREREQzMzNEREREREREREREREREREREREREREREREQzMzNEREREREREREREREQzMzMzMzMiIiIzMzMzMzMzMzMzMzNERERERERERERVVVVVVVVVVVVmZmZ3d3eqqqq7u7u7u7vd3d3///////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3dzMzM3d3d7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d7u7u3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3dzMzMu7u7qqqqqqqqmZmZmZmZmZmZiIiIiIiIiIiId3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3ZmZmd3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVZmZmd3d3ZmZmd3d3d3d3ZmZmd3d3iIiId3d3d3d3iIiId3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3iIiId3d3iIiId3d3iIiId3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREVVVVREREREREREREREREREREREREREREREREREREMzMzREREVVVVVVVVZmZmZmZmZmZmVVVVVVVVd3d3iIiIiIiId3d3d3d3VVVVZmZmd3d3iIiId3d3ZmZmVVVVREREVVVVd3d3iIiId3d3ZmZmVVVVZmZmZmZmiIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3VVVVVVVVVVVVVVVVREREMzMzREREREREVVVVmZmZzMzMqqqqiIiId3d3iIiImZmZu7u73d3dzMzMzMzMu7u7qqqqqqqqqqqqqqqqzMzM3d3dzMzMzMzMu7u7zMzMzMzMu7u7mZmZmZmZqqqqqqqqiIiIiIiImZmZmZmZqqqqqqqqqqqqmZmZmZmZqqqqqqqqiIiIZmZmVVVVREREREREVVVVmZmZqqqqqqqqqqqqqqqqu7u7u7u7u7u7qqqqqqqqqqqqu7u7zMzMzMzMu7u7mZmZiIiIiIiImZmZu7u7zMzMzMzMu7u7u7u7u7u7zMzMu7u7u7u73d3du7u7qqqqqqqqqqqqu7u7u7u7mZmZd3d3mZmZzMzMzMzMzMzMu7u7qqqqqqqqmZmZiIiImZmZmZmZmZmZmZmZmZmZmZmZiIiIZmZmZmZmiIiIqqqqzMzMzMzMzMzMqqqqqqqqmZmZmZmZmZmZiIiId3d3ZmZmd3d3iIiId3d3VVVVREREVVVViIiIu7u7mZmZmZmZmZmZqqqqqqqqqqqqmZmZmZmZiIiIZmZmd3d3ZmZmZmZmREREREREmZmZzMzMzMzMu7u7mZmZu7u7qqqqqqqqqqqqqqqqmZmZmZmZmZmZiIiIiIiId3d3d3d3ZmZmiIiIqqqqqqqqmZmZmZmZmZmZmZmZmZmZd3d3mZmZiIiId3d3ZmZmZmZmZmZmVVVVREREZmZmiIiImZmZiIiIiIiImZmZiIiId3d3d3d3mZmZqqqqqqqqu7u7qqqqqqqqmZmZmZmZmZmZqqqqmZmZmZmZmZmZmZmZmZmZd3d3d3d3ZmZmd3d3iIiIiIiId3d3d3d3d3d3iIiId3d3d3d3ZmZmVVVVZmZmZmZmVVVVZmZmVVVVMzMzMzMzMzMzREREREREREREREREVVVVd3d3iIiId3d3iIiImZmZu7u7qqqqqqqqd3d3ZmZmZmZmZmZmVVVVZmZmd3d3d3d3ZmZmd3d3d3d3iIiIZmZmZmZmZmZmd3d3iIiIqqqqmZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3d3d3iIiId3d3ZmZmd3d3ZmZmVVVVZmZmd3d3mZmZmZmZiIiId3d3ZmZmVVVVREREREREVVVVVVVVZmZmZmZmZmZmZmZmd3d3ZmZmZmZmREREREREMzMzMzMzVVVVmZmZqqqqiIiId3d3ZmZmVVVVREREREREZmZmZmZmZmZmZmZmREREVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVd3d3d3d3d3d3ZmZmREREREREREREVVVVVVVVVVVVVVVVZmZmZmZmVVVVREREVVVVVVVVVVVVREREREREREREREREVVVVZmZmVVVVREREREREVVVVREREREREREREVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzREREVVVVVVVVREREREREREREREREREREREREZmZmVVVVREREREREREREREREMzMzMzMzMzMzMzMzREREREREREREMzMzREREVVVVVVVVREREREREREREREREMzMzREREd3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVVVVVREREREREMzMzREREREREREREVVVVVVVVREREREREMzMzREREREREREREREREMzMzREREMzMzIiIiIiIiMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzREREREREVVVVREREVVVVREREMzMzMzMzREREVVVVREREVVVVREREREREREREREREREREREREREREREREMzMzREREREREVVVVVVVVVVVVREREREREREREREREMzMzREREZmZmVVVVREREREREREREVVVVREREREREREREREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzZmZmZmZmREREMzMzREREREREMzMzREREVVVVVVVVZmZmREREREREMzMzREREREREREREZmZmqqqqd3d3REREREREREREREREREREREREREREREREREREZmZmZmZmZmZmd3d3ZmZmVVVVIiIiMzMzMzMzMzMzZmZmd3d3qqqqqqqqd3d3VVVVZmZmZmZmREREIiIiIiIiIiIiIiIiIiIiMzMzMzMzVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVREREREREVVVVREREVVVVREREREREMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVREREVVVVREREREREREREREREVVVVREREREREREREREREVVVVREREREREVVVVVVVVVVVVZmZmZmZmZmZmVVVVREREREREVVVVREREREREREREREREd3d3ZmZmREREREREVVVVZmZmZmZmZmZmZmZmVVVViIiIqqqqiIiIREREIiIiVVVVu7u7u7u7d3d3ZmZmZmZmVVVVZmZmVVVVREREVVVVREREREREREREMzMzREREVVVVVVVVREREREREVVVVREREVVVVd3d3d3d3d3d3iIiIiIiImZmZiIiId3d3ZmZmVVVVVVVVREREREREVVVVZmZmd3d3d3d3iIiIqqqqiIiId3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiId3d3ZmZmZmZmd3d3ZmZmVVVVVVVVREREREREVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmVVVVZmZmd3d3iIiIu7u7zMzMu7u7mZmZiIiId3d3d3d3ZmZmZmZmd3d3d3d3d3d3d3d3ZmZmZmZmd3d3ZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVZmZmZmZmVVVVVVVVVVVVREREVVVVVVVViIiIiIiId3d3d3d3iIiIiIiId3d3iIiId3d3mZmZu7u7zMzMqqqqiIiIiIiId3d3mZmZu7u7u7u7d3d3ZmZmZmZmZmZmVVVVZmZmd3d3d3d3d3d3mZmZd3d3VVVVVVVVREREREREMzMzMzMzMzMzMzMzVVVVREREREREREREREREREREREREREREMzMzIiIiIiIiMzMzMzMzMzMzMzMzREREREREREREREREREREVVVVZmZmZmZmiIiIu7u7u7u7zMzM7u7u////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7t3d3czMzN3d3e7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3d3d3e7u7t3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3czMzMzMzKqqqpmZmYiIiHd3d3d3d2ZmZlVVVWZmZlVVVVVVVWZmZmZmZmZmZlVVVURERERERFVVVURERERERERERFVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiJmZmYiIiJmZmYiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZkRERFVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVURERERERFVVVWZmZmZmZlVVVVVVVVVVVVVVVXd3d3d3d2ZmZmZmZmZmZlVVVVVVVYiIiIiIiGZmZlVVVWZmZmZmZlVVVXd3d3d3d4iIiHd3d3d3d3d3d3d3d2ZmZlVVVVVVVVVVVURERERERFVVVURERERERFVVVZmZmbu7u6qqqmZmZmZmZpmZmbu7u8zMzLu7u8zMzMzMzLu7u6qqqqqqqqqqqqqqqszMzMzMzN3d3bu7u7u7u8zMzLu7u6qqqpmZmaqqqqqqqpmZmZmZmZmZmZmZmaqqqqqqqpmZmZmZmYiIiKqqqqqqqoiIiHd3d2ZmZlVVVVVVVURERHd3d6qqqqqqqpmZmaqqqqqqqru7u7u7u7u7u6qqqpmZmaqqqru7u8zMzLu7u7u7u6qqqpmZmaqqqpmZmczMzMzMzMzMzLu7u7u7u7u7u8zMzMzMzMzMzMzMzLu7u6qqqru7u6qqqqqqqqqqqpmZmXd3d7u7u8zMzMzMzLu7u7u7u7u7u6qqqoiIiHd3d4iIiIiIiIiIiIiIiHd3d4iIiIiIiHd3d3d3d3d3d7u7u8zMzMzMzLu7u5mZmZmZmZmZmYiIiJmZmYiIiJmZmWZmZnd3d4iIiGZmZlVVVURERERERIiIiKqqqru7u6qqqpmZmZmZmZmZmYiIiJmZmZmZmYiIiHd3d2ZmZmZmZlVVVURERFVVVZmZmczMzMzMzMzMzKqqqqqqqqqqqpmZmaqqqru7u6qqqpmZmZmZmYiIiHd3d2ZmZmZmZmZmZnd3d5mZmZmZmYiIiHd3d4iIiJmZmXd3d3d3d4iIiHd3d2ZmZmZmZnd3d1VVVURERFVVVWZmZmZmZoiIiIiIiHd3d3d3d2ZmZnd3d5mZmaqqqru7u7u7u8zMzKqqqqqqqpmZmZmZmaqqqpmZmZmZmZmZmZmZmaqqqpmZmYiIiGZmZmZmZnd3d5mZmXd3d3d3d4iIiIiIiHd3d2ZmZlVVVVVVVWZmZpmZmYiIiFVVVVVVVVVVVURERDMzMzMzM0RERERERFVVVVVVVVVVVXd3d3d3d3d3d4iIiKqqqru7u6qqqoiIiHd3d2ZmZmZmZmZmZlVVVWZmZnd3d4iIiGZmZnd3d4iIiIiIiFVVVWZmZmZmZmZmZpmZmaqqqqqqqoiIiJmZmYiIiHd3d4iIiIiIiHd3d4iIiHd3d3d3d4iIiIiIiIiIiHd3d3d3d4iIiGZmZlVVVWZmZnd3d4iIiJmZmZmZmWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d2ZmZlVVVTMzMzMzMzMzMzMzM2ZmZoiIiJmZmYiIiGZmZmZmZlVVVURERERERFVVVVVVVWZmZlVVVVVVVURERFVVVWZmZmZmZmZmZlVVVVVVVVVVVURERFVVVXd3d3d3d2ZmZmZmZkRERFVVVURERERERFVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVURERERERFVVVURERDMzM0RERGZmZmZmZlVVVVVVVURERERERERERFVVVURERERERERERFVVVURERERERFVVVWZmZlVVVVVVVURERFVVVVVVVURERERERFVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERERERERERDMzM0RERERERERERERERERERERERERERFVVVURERDMzMzMzMzMzMyIiIjMzM0RERERERERERERERDMzM0RERFVVVVVVVURERERERERERERERDMzM0RERGZmZmZmZlVVVVVVVURERERERERERERERERERDMzM0RERFVVVVVVVVVVVURERDMzM0RERERERDMzM0RERGZmZlVVVVVVVURERERERDMzM0RERERERERERDMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzM0RERERERERERERERERERERERERERERERDMzM0RERERERERERERERFVVVURERFVVVURERERERERERDMzM0RERDMzM0RERERERFVVVVVVVURERERERERERDMzMzMzMzMzM0RERFVVVURERDMzM0RERFVVVVVVVURERERERDMzM0RERFVVVURERERERERERERERDMzMzMzMzMzMzMzMzMzM1VVVXd3d0RERERERERERERERERERERERERERGZmZlVVVURERERERDMzMzMzM0RERERERGZmZqqqqoiIiFVVVURERFVVVVVVVURERFVVVURERFVVVVVVVVVVVXd3d3d3d3d3d3d3d1VVVTMzMyIiIjMzMzMzM1VVVYiIiIiIiIiIiHd3d1VVVVVVVXd3d1VVVTMzMyIiIiIiIiIiIhERETMzM0RERERERFVVVWZmZlVVVVVVVVVVVWZmZmZmZmZmZlVVVURERFVVVVVVVVVVVURERERERERERERERFVVVVVVVURERERERDMzMyIiIjMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERFVVVVVVVURERERERERERERERERERERERERERERERERERERERERERERERFVVVVVVVVVVVWZmZlVVVVVVVURERERERERERERERFVVVVVVVURERFVVVXd3d2ZmZlVVVVVVVVVVVWZmZmZmZnd3d3d3d2ZmZoiIiKqqqoiIiERERDMzM1VVVbu7u8zMzHd3d2ZmZlVVVVVVVWZmZlVVVVVVVURERERERFVVVURERERERERERERERFVVVVVVVURERFVVVURERFVVVXd3d4iIiJmZmYiIiIiIiIiIiIiIiIiIiFVVVVVVVVVVVVVVVVVVVURERFVVVVVVVXd3d4iIiIiIiIiIiIiIiGZmZnd3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVURERERERFVVVWZmZlVVVWZmZnd3d2ZmZmZmZoiIiJmZmYiIiKqqqszMzLu7u5mZmZmZmXd3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d2ZmZmZmZmZmZlVVVVVVVURERFVVVVVVVURERFVVVWZmZkRERGZmZlVVVVVVVURERFVVVWZmZoiIiIiIiHd3d2ZmZnd3d4iIiKqqqqqqqqqqqru7u6qqqqqqqoiIiHd3d3d3d5mZmbu7u6qqqnd3d2ZmZmZmZlVVVVVVVVVVVWZmZmZmZoiIiLu7u4iIiFVVVWZmZlVVVURERDMzM0RERDMzM0RERERERERERERERERERERERDMzM0RERDMzMzMzMyIiIjMzMyIiIjMzMzMzM0RERERERERERFVVVVVVVURERFVVVWZmZmZmZoiIiKqqqszMzP///////+7u7v///////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7d3d3d3d3d3d3u7u7u7u7u7u7d3d3u7u7d3d3u7u7d3d3u7u7d3d3u7u7d3d3u7u7d3d3d3d3MzMzMzMy7u7uqqqq7u7uqqqq7u7vMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzd3d3MzMzMzMzMzMy7u7u7u7uZmZmZmZl3d3dmZmZmZmZmZmZVVVVVVVVmZmZVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVERERVVVVERERVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3dmZmZmZmZ3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIh3d3eIiIh3d3d3d3d3d3eIiIh3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3dmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVERERERERVVVVmZmZmZmZVVVVERERERERERERERERERERVVVVVVVVVVVVVVVWIiIiIiIh3d3dmZmZ3d3eIiIhVVVVmZmZ3d3eIiIiIiIh3d3d3d3dmZmZmZmZmZmZVVVVERERERERERERVVVVVVVVERERVVVWZmZm7u7uZmZlmZmZmZmaqqqrMzMzMzMy7u7vMzMzMzMy7u7uqqqqqqqqqqqqqqqq7u7vMzMzMzMzMzMzMzMzMzMy7u7uqqqq7u7u7u7uqqqqqqqqIiIiZmZmqqqq7u7uZmZmZmZmZmZmIiIiZmZmqqqqIiIiIiIh3d3dVVVVERERVVVWZmZm7u7uqqqqqqqqqqqq7u7u7u7u7u7uqqqqqqqqZmZm7u7u7u7u7u7vMzMzMzMyqqqqZmZmIiIiZmZnMzMzd3d3MzMzMzMy7u7vMzMzMzMzMzMy7u7u7u7uZmZmqqqq7u7u7u7uqqqqZmZmZmZmIiIi7u7vMzMzMzMy7u7uqqqrMzMyqqqqIiIh3d3eIiIiIiIiIiIh3d3d3d3eIiIiZmZl3d3dmZmZ3d3eZmZnMzMy7u7u7u7uZmZmIiIiIiIiZmZm7u7uZmZmIiIh3d3d3d3eIiIh3d3dVVVVVVVVERERmZmaqqqrMzMyqqqqZmZmIiIiIiIiIiIh3d3d3d3eIiIiIiIhmZmZVVVVVVVVVVVVERER3d3e7u7vd3d27u7uqqqqqqqp3d3eIiIiqqqqqqqqZmZmZmZmZmZl3d3d3d3dmZmZVVVVERER3d3eIiIiZmZmIiIh3d3d3d3eIiIiIiIh3d3eIiIh3d3d3d3d3d3d3d3dVVVVERERERERVVVV3d3d3d3d3d3d3d3dmZmZ3d3eIiIiIiIiqqqq7u7vMzMy7u7uqqqqqqqqZmZmqqqqqqqqZmZmIiIiqqqq7u7uqqqqZmZl3d3dmZmZmZmZ3d3eIiIiIiIh3d3d3d3d3d3eIiIhmZmZVVVVERERmZmaZmZl3d3dmZmZmZmZVVVVEREQzMzMzMzNERERERERVVVVVVVV3d3d3d3dmZmZ3d3eIiIiZmZm7u7uqqqqZmZlmZmZmZmZmZmZVVVVVVVV3d3eIiIh3d3d3d3d3d3d3d3eIiIhmZmZmZmZVVVVmZmaZmZmqqqqqqqqZmZmIiIiIiIiIiIiIiIh3d3eIiIiIiIh3d3d3d3eIiIiIiIh3d3d3d3eIiIiIiIhmZmZVVVVmZmZ3d3eqqqqqqqqIiIhmZmZVVVVERERVVVVVVVVVVVVVVVVVVVV3d3dmZmZ3d3dmZmZEREREREQzMzMzMzMzMzMzMzNVVVVVVVVmZmZ3d3d3d3d3d3dERERERERERERERERERERERERVVVVERERVVVVERER3d3eIiIhmZmZmZmZVVVVVVVVEREQzMzN3d3d3d3dmZmZVVVVmZmZVVVVERERERERERERVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERERERmZmZVVVVVVVVEREREREREREREREREREREREREREREREQzMzNVVVVmZmZmZmZERERERERVVVVVVVVEREREREREREREREREREREREQzMzNEREQzMzMzMzNEREQzMzNEREREREREREQzMzNERERERERVVVVEREREREREREREREREREREREQzMzMzMzMzMzNEREREREREREQzMzMiIiIzMzMiIiIiIiIzMzMzMzNEREQzMzMzMzNERERVVVVEREQzMzNEREREREQzMzNERERERERVVVVVVVVVVVVVVVVEREREREREREQzMzNEREREREREREREREREREQzMzMzMzNERERERERERERERERVVVVVVVVEREREREREREREREREREREREQzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzMzMzNEREREREREREREREREREREREQzMzNERERERERERERERERERERERERERERVVVVEREREREREREREREREREQzMzNERERERERVVVVVVVVERERVVVVERERVVVVEREQzMzNEREREREREREQzMzNERERERERVVVVERERERERERERERERERERVVVVVVVVVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzNERER3d3dVVVVERERVVVVVVVVVVVVERERERERVVVVVVVVEREREREQzMzMzMzMzMzNERERmZmaZmZmIiIhmZmZERERVVVVVVVVVVVVERERERERERERVVVVmZmZ3d3d3d3d3d3eIiIhmZmYzMzMzMzMzMzMzMzNERER3d3d3d3d3d3d3d3dmZmZVVVVmZmZ3d3dVVVUzMzMREREiIiIiIiIiIiJERERERERVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZVVVVmZmZVVVVVVVVVVVVERERERERERERERERERERVVVVEREREREQzMzMzMzMzMzMzMzNEREREREQzMzNEREREREQzMzNEREQzMzMzMzNERERERERERERERERERERERERVVVVEREQzMzNERERVVVVERERVVVVERERERERVVVVERERVVVVVVVVVVVVVVVVmZmZVVVVEREQzMzNERERERERERERERERERERERERVVVVmZmZmZmZmZmZERERVVVVmZmZ3d3d3d3d3d3d3d3eqqqq7u7uIiIhVVVUiIiJVVVW7u7vMzMyIiIhVVVVmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVEREQzMzNVVVVVVVVVVVVERERERERERERVVVVVVVVmZmaIiIiZmZmZmZl3d3d3d3d3d3d3d3dmZmZVVVVVVVVVVVVERERVVVVERERVVVVVVVVmZmZmZmZmZmZ3d3d3d3d3d3d3d3eIiIh3d3d3d3eIiIiIiIiIiIiIiIh3d3eIiIhmZmZmZmZmZmZmZmZ3d3dmZmZVVVVmZmZ3d3d3d3d3d3eIiIh3d3d3d3eIiIiIiIiIiIiIiIiZmZmZmZmZmZmZmZmIiIh3d3d3d3d3d3dmZmZ3d3eIiIiZmZmZmZl3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERERERmZmZmZmZ3d3dmZmZmZmZ3d3eqqqqqqqq7u7uqqqq7u7uqqqqZmZmIiIhmZmZ3d3eIiIiqqqqZmZl3d3dmZmZVVVVVVVVVVVVERERVVVV3d3eqqqq7u7uZmZl3d3eIiIhmZmZEREREREREREREREREREREREREREREREREREREREREREQzMzMiIiIiIiIzMzMiIiIzMzMzMzMzMzNEREQzMzNERERERERVVVVVVVVVVVVVVVVmZmaZmZmqqqrd3d3///////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////7u7u3d3dzMzMu7u7zMzM3d3d3d3d7u7u3d3d3d3d3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMu7u7u7u7qqqqqqqqu7u7u7u7zMzMzMzMzMzM3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzM3d3dzMzMzMzM3d3dzMzMzMzMu7u7u7u7qqqqqqqqqqqqqqqqqqqqmZmZqqqqqqqqqqqqmZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZmZmZmZmZqqqqmZmZiIiIiIiIiIiIiIiId3d3mZmZiIiIiIiImZmZiIiImZmZiIiImZmZiIiIiIiIiIiIiIiIiIiId3d3iIiId3d3d3d3d3d3d3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3iIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3iIiIiIiId3d3d3d3d3d3iIiIiIiIiIiId3d3d3d3iIiId3d3d3d3ZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiId3d3iIiId3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3d3d3ZmZmd3d3ZmZmd3d3ZmZmVVVVZmZmd3d3ZmZmVVVVVVVVREREREREVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmd3d3iIiIiIiId3d3ZmZmVVVVZmZmiIiId3d3ZmZmZmZmVVVVREREVVVVVVVVREREREREREREREREREREVVVVVVVVd3d3u7u7qqqqd3d3ZmZmu7u7zMzMzMzMu7u7zMzMzMzMzMzMu7u7qqqqqqqqmZmZqqqqu7u7qqqqu7u73d3dzMzMqqqqu7u7zMzMu7u7qqqqmZmZiIiIiIiImZmZmZmZiIiIiIiIiIiIqqqqqqqqiIiId3d3d3d3d3d3VVVVVVVVd3d3u7u7zMzMmZmZmZmZqqqqu7u7u7u7zMzMu7u7u7u7u7u7qqqqu7u7mZmZqqqqzMzMzMzMiIiIZmZmmZmZ3d3dzMzMzMzMzMzMzMzMzMzMzMzM3d3du7u7qqqqqqqqu7u7u7u7u7u7qqqqiIiId3d3iIiIu7u7zMzM3d3du7u7qqqqqqqqmZmZiIiImZmZiIiImZmZmZmZiIiId3d3iIiId3d3d3d3ZmZmZmZmZmZmmZmZqqqqqqqqiIiImZmZd3d3iIiIqqqqmZmZd3d3ZmZmd3d3ZmZmVVVVZmZmVVVVREREVVVViIiIqqqqmZmZiIiIiIiIiIiId3d3d3d3iIiImZmZd3d3ZmZmVVVVZmZmZmZmREREVVVViIiIqqqqmZmZiIiIiIiId3d3iIiIiIiIiIiIiIiIiIiImZmZiIiId3d3VVVVREREVVVVd3d3iIiIiIiId3d3d3d3d3d3iIiId3d3iIiId3d3d3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVZmZmiIiIiIiId3d3d3d3d3d3d3d3mZmZqqqqu7u7u7u7u7u7qqqqmZmZiIiIqqqqqqqqmZmZmZmZqqqqmZmZd3d3ZmZmd3d3ZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3VVVVREREVVVVd3d3d3d3VVVVZmZmZmZmVVVVMzMzREREREREREREREREREREZmZmd3d3ZmZmZmZmiIiIiIiIiIiIqqqqqqqqmZmZiIiId3d3ZmZmVVVVVVVVZmZmZmZmVVVVZmZmd3d3mZmZd3d3d3d3iIiIZmZmZmZmd3d3mZmZu7u7qqqqmZmZiIiId3d3ZmZmd3d3d3d3iIiIiIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3ZmZmd3d3mZmZmZmZd3d3ZmZmZmZmREREVVVVREREREREVVVVZmZmZmZmd3d3ZmZmVVVVREREMzMzMzMzREREREREREREMzMzMzMzREREd3d3d3d3VVVVREREREREVVVVREREREREVVVVVVVVVVVVREREVVVVZmZmZmZmZmZmVVVVVVVVMzMzREREREREZmZmZmZmZmZmVVVVVVVVREREREREREREVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVREREREREREREMzMzMzMzREREVVVVREREREREVVVVREREREREREREMzMzREREMzMzREREREREREREVVVVZmZmVVVVREREVVVVVVVVREREMzMzMzMzMzMzREREREREREREREREVVVVVVVVMzMzMzMzREREREREMzMzREREREREREREVVVVVVVVVVVVREREMzMzREREMzMzMzMzIiIiMzMzREREMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzREREREREVVVVREREMzMzREREREREREREMzMzREREREREVVVVVVVVVVVVREREMzMzMzMzMzMzMzMzREREVVVVREREMzMzMzMzREREREREREREREREREREVVVVVVVVREREREREREREREREMzMzREREMzMzMzMzMzMzREREMzMzMzMzIiIiMzMzMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiMzMzREREVVVVREREVVVVVVVVREREREREMzMzREREMzMzREREMzMzMzMzREREVVVVREREREREVVVVREREREREREREREREVVVVVVVVVVVVREREREREREREREREREREREREMzMzMzMzMzMzREREREREVVVVVVVVREREREREREREREREVVVVVVVVVVVVVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzZmZmZmZmVVVVVVVVMzMzREREREREREREZmZmZmZmREREREREREREREREMzMzMzMzZmZmiIiIZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVREREZmZmZmZmd3d3iIiIZmZmREREIiIiMzMzMzMzZmZmd3d3iIiIiIiId3d3ZmZmVVVVVVVVd3d3ZmZmREREMzMzIiIiIiIiIiIiMzMzREREVVVVVVVVZmZmd3d3d3d3ZmZmZmZmZmZmd3d3ZmZmZmZmVVVVVVVVVVVVREREREREREREVVVVVVVVREREREREREREREREMzMzMzMzREREREREREREREREMzMzREREMzMzMzMzREREREREREREREREREREREREREREREREVVVVREREMzMzREREVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVMzMzMzMzREREREREREREVVVVVVVVREREREREVVVVZmZmVVVVZmZmVVVVVVVVd3d3iIiImZmZd3d3iIiIzMzMzMzMmZmZVVVVIiIiVVVVqqqqu7u7d3d3ZmZmVVVVVVVVVVVVZmZmVVVVREREREREVVVVREREVVVVVVVVVVVVREREREREVVVVREREVVVVVVVVZmZmiIiIiIiIiIiId3d3VVVVZmZmd3d3VVVVVVVVZmZmZmZmVVVVVVVVREREVVVVREREVVVVVVVVZmZmZmZmZmZmZmZmd3d3ZmZmd3d3d3d3d3d3mZmZmZmZiIiIiIiIiIiIiIiId3d3ZmZmZmZmd3d3ZmZmZmZmZmZmd3d3iIiImZmZmZmZmZmZqqqqmZmZiIiId3d3d3d3d3d3d3d3iIiIiIiIiIiId3d3d3d3d3d3d3d3ZmZmd3d3iIiIiIiImZmZd3d3ZmZmZmZmZmZmVVVVVVVVREREREREREREVVVVZmZmVVVVVVVVVVVVREREREREREREREREZmZmVVVVZmZmd3d3mZmZqqqqu7u7mZmZqqqqu7u7qqqqmZmZiIiIZmZmZmZmd3d3iIiIqqqqd3d3VVVVREREREREREREVVVVZmZmqqqq7u7u3d3dqqqqmZmZiIiId3d3ZmZmVVVVREREVVVVREREREREREREREREREREREREREREIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREVVVVVVVVZmZmZmZmd3d3qqqq3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7t3d3czMzLu7u7u7u8zMzN3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3e7u7t3d3d3d3d3d3e7u7t3d3e7u7t3d3d3d3czMzMzMzN3d3czMzN3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3d3d3d3d3e7u7u7u7u7u7t3d3d3d3d3d3czMzMzMzMzMzLu7u7u7u6qqqqqqqqqqqqqqqpmZmYiIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiJmZmZmZmZmZmZmZmaqqqqqqqpmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiJmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiIiIiJmZmYiIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d4iIiHd3d4iIiIiIiHd3d4iIiIiIiIiIiHd3d4iIiIiIiIiIiIiIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiHd3d3d3d3d3d4iIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZnd3d3d3d2ZmZnd3d3d3d3d3d4iIiHd3d3d3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d3d3d2ZmZmZmZlVVVVVVVVVVVURERERERGZmZmZmZlVVVWZmZlVVVURERFVVVXd3d4iIiIiIiGZmZnd3d2ZmZmZmZnd3d3d3d2ZmZnd3d1VVVURERDMzM0RERFVVVVVVVVVVVURERFVVVURERERERGZmZpmZmaqqqnd3d3d3d8zMzMzMzLu7u7u7u8zMzLu7u8zMzKqqqqqqqpmZmYiIiHd3d5mZmbu7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqqqqqpmZmZmZmYiIiIiIiHd3d3d3d4iIiJmZmbu7u5mZmYiIiHd3d2ZmZlVVVVVVVWZmZnd3d7u7u8zMzLu7u6qqqoiIiJmZmaqqqru7u6qqqru7u7u7u6qqqqqqqpmZmYiIiKqqqqqqqnd3d2ZmZoiIiN3d3czMzMzMzMzMzLu7u8zMzN3d3bu7u7u7u6qqqqqqqqqqqqqqqqqqqpmZmWZmZmZmZmZmZoiIiLu7u93d3bu7u6qqqpmZmYiIiJmZmaqqqpmZmaqqqqqqqoiIiIiIiIiIiHd3d2ZmZmZmZlVVVVVVVYiIiIiIiIiIiHd3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiHd3d2ZmZlVVVWZmZkRERFVVVWZmZnd3d3d3d3d3d3d3d4iIiIiIiIiIiJmZmZmZmYiIiIiIiIiIiIiIiHd3d1VVVURERFVVVYiIiJmZmYiIiIiIiJmZmYiIiIiIiJmZmYiIiIiIiIiIiHd3d3d3d1VVVVVVVWZmZnd3d3d3d6qqqpmZmYiIiHd3d3d3d2ZmZoiIiIiIiHd3d3d3d3d3d1VVVVVVVWZmZlVVVXd3d5mZmZmZmZmZmZmZmZmZmYiIiIiIiKqqqqqqqru7u7u7u6qqqpmZmZmZmYiIiJmZmaqqqqqqqqqqqpmZmXd3d3d3d2ZmZmZmZmZmZnd3d2ZmZnd3d4iIiHd3d3d3d3d3d2ZmZlVVVURERERERHd3d3d3d1VVVVVVVURERFVVVURERERERERERFVVVURERFVVVVVVVWZmZmZmZmZmZoiIiIiIiGZmZpmZmaqqqqqqqoiIiHd3d1VVVVVVVURERFVVVVVVVVVVVWZmZoiIiIiIiHd3d5mZmZmZmWZmZlVVVVVVVXd3d6qqqqqqqoiIiHd3d2ZmZmZmZmZmZnd3d4iIiIiIiIiIiIiIiHd3d4iIiHd3d4iIiHd3d4iIiHd3d2ZmZmZmZnd3d4iIiHd3d3d3d1VVVVVVVURERERERERERFVVVXd3d2ZmZmZmZlVVVURERDMzM0RERERERERERDMzMzMzMzMzMyIiIjMzM2ZmZnd3d2ZmZlVVVVVVVURERERERFVVVVVVVVVVVURERFVVVWZmZnd3d2ZmZmZmZmZmZlVVVTMzM0RERFVVVVVVVWZmZmZmZmZmZlVVVVVVVURERDMzM0RERFVVVVVVVVVVVWZmZmZmZkRERFVVVURERDMzM0RERDMzM0RERERERERERERERFVVVURERFVVVURERERERERERDMzM0RERDMzM0RERERERGZmZlVVVURERERERFVVVWZmZkRERDMzMzMzMzMzM0RERERERERERERERFVVVURERDMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVVVVVURERERERERERDMzMzMzMyIiIjMzMzMzM0RERDMzM0RERERERDMzMzMzMyIiIjMzMzMzMzMzMyIiIiIiIjMzMzMzM0RERFVVVURERERERERERERERERERDMzM0RERERERERERERERFVVVURERERERERERDMzM0RERDMzM0RERERERDMzMzMzM0RERFVVVURERFVVVVVVVURERERERERERERERDMzM0RERDMzM0RERDMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIhERETMzMzMzM0RERERERERERERERFVVVURERERERDMzMzMzM0RERDMzMzMzMzMzMzMzM0RERERERERERERERERERERERERERFVVVVVVVVVVVURERFVVVURERERERERERERERDMzMzMzM0RERDMzMzMzM0RERERERFVVVURERERERERERERERFVVVVVVVVVVVVVVVURERERERERERDMzMzMzMzMzMzMzMzMzMzMzM0RERGZmZkRERERERDMzMzMzM0RERERERGZmZnd3d1VVVTMzM0RERFVVVTMzMzMzM1VVVYiIiIiIiFVVVWZmZlVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVVVVVWZmZnd3d1VVVURERCIiIjMzM0RERIiIiHd3d3d3d3d3d3d3d2ZmZmZmZkRERERERFVVVVVVVTMzMzMzMyIiIiIiIjMzMzMzM0RERGZmZnd3d4iIiIiIiHd3d2ZmZmZmZnd3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERDMzM0RERERERERERERERERERERERDMzMzMzM0RERDMzM0RERERERERERERERFVVVVVVVVVVVURERERERFVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVTMzMzMzM0RERERERERERFVVVURERFVVVVVVVURERFVVVVVVVWZmZlVVVVVVVXd3d3d3d6qqqpmZmXd3d4iIiMzMzMzMzJmZmVVVVTMzM0RERJmZmaqqqmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVURERERERERERFVVVVVVVURERFVVVURERFVVVURERFVVVVVVVWZmZmZmZnd3d3d3d2ZmZmZmZmZmZnd3d2ZmZlVVVVVVVWZmZlVVVWZmZlVVVURERERERERERERERFVVVWZmZmZmZmZmZnd3d2ZmZnd3d3d3d3d3d4iIiIiIiIiIiHd3d4iIiIiIiGZmZlVVVXd3d3d3d3d3d3d3d3d3d3d3d4iIiJmZmYiIiIiIiIiIiJmZmZmZmYiIiGZmZmZmZnd3d3d3d4iIiIiIiHd3d3d3d3d3d1VVVURERERERGZmZpmZmczMzJmZmXd3d2ZmZlVVVVVVVURERDMzM0RERERERERERERERGZmZmZmZlVVVURERERERFVVVVVVVVVVVWZmZmZmZmZmZpmZmaqqqpmZmZmZmaqqqszMzLu7u5mZmXd3d2ZmZlVVVWZmZnd3d4iIiHd3d1VVVVVVVURERFVVVXd3d3d3d8zMzN3d3d3d3czMzJmZmYiIiHd3d3d3d3d3d3d3d1VVVVVVVVVVVVVVVURERERERDMzMzMzMyIiIiIiIiIiIjMzM0RERDMzMzMzM0RERDMzM0RERERERERERERERFVVVWZmZnd3d4iIiKqqqt3d3f///////////////////+7u7v///////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3u7u7d3d3d3d3u7u7d3d3d3d3u7u7d3d3u7u7d3d3u7u7d3d3u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMyqqqqqqqqqqqqZmZmIiIiIiIh3d3d3d3dmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiZmZm7u7uqqqqIiIiZmZmZmZmIiIiZmZmIiIiIiIiZmZmZmZmZmZmIiIiZmZmIiIiZmZmIiIiIiIiIiIh3d3d3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3dmZmZ3d3dmZmZ3d3dmZmZ3d3d3d3dmZmZ3d3dmZmZ3d3d3d3d3d3d3d3dmZmZ3d3d3d3dmZmZmZmZ3d3d3d3dmZmZ3d3dmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZVVVVVVVVERERVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZVVVV3d3dmZmZmZmZmZmZVVVVVVVVVVVVmZmZVVVVmZmZVVVVVVVVERER3d3eIiIh3d3dmZmZ3d3d3d3d3d3dmZmZmZmZ3d3d3d3dVVVUzMzNERERVVVVmZmZmZmZERERVVVVERERVVVVERERVVVWIiIi7u7t3d3eZmZnd3d3MzMy7u7uqqqqqqqq7u7u7u7uqqqqqqqqZmZmZmZmIiIiIiIiqqqqqqqqZmZmZmZm7u7vMzMy7u7uqqqqZmZmZmZmZmZmZmZl3d3d3d3d3d3eZmZmZmZmqqqqZmZmIiIh3d3dmZmZERERERERERER3d3e7u7vMzMy7u7u7u7uqqqqZmZmZmZmqqqqZmZmZmZmIiIiZmZmZmZmqqqqIiIiIiIiIiIhmZmZVVVWIiIi7u7u7u7u7u7u7u7u7u7u7u7vMzMzMzMyqqqqqqqq7u7uqqqqqqqqZmZmIiIhmZmZVVVVERERmZmaZmZmqqqq7u7uqqqqqqqqIiIiqqqq7u7u7u7vMzMyqqqqqqqqZmZmIiIiIiIhmZmZERERVVVV3d3eZmZmZmZmIiIhmZmZmZmZmZmZ3d3eZmZmZmZmZmZmZmZmZmZmIiIiIiIhVVVVVVVVERERVVVVVVVVmZmZmZmZ3d3dmZmZ3d3d3d3eZmZmqqqqZmZmIiIiIiIiIiIiZmZmZmZlVVVVERERmZmaIiIiIiIiIiIiIiIiIiIiIiIiZmZmZmZmZmZmIiIiIiIh3d3dmZmZmZmZVVVWIiIiIiIiqqqqqqqqZmZmIiIiIiIh3d3d3d3eIiIiZmZl3d3eIiIh3d3dmZmZVVVVmZmZmZmZ3d3eZmZm7u7uZmZmqqqqZmZmZmZmZmZmqqqqZmZmqqqq7u7u7u7uqqqqqqqqqqqqqqqq7u7uZmZmIiIh3d3dmZmZ3d3d3d3d3d3eIiIh3d3d3d3eIiIiIiIiIiIiIiIh3d3dmZmZVVVVVVVVERER3d3dmZmZVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVERERVVVVmZmZmZmZ3d3eZmZl3d3dmZmZ3d3eqqqqqqqqIiIhmZmZVVVVERERVVVVVVVVVVVVmZmZ3d3eZmZl3d3eIiIiqqqp3d3d3d3dmZmZmZmZ3d3eZmZmqqqqZmZmIiIh3d3dmZmZVVVVmZmZ3d3eIiIiIiIh3d3eIiIh3d3eIiIiZmZmZmZmIiIh3d3dmZmZmZmaIiIiZmZl3d3dmZmZVVVVVVVVERERERERERERERERVVVVmZmZVVVVVVVVVVVVEREREREREREREREREREQzMzMzMzMzMzMzMzNERERmZmZ3d3dmZmZEREREREREREQzMzNERERERERERERmZmZ3d3dmZmZmZmZmZmZ3d3dVVVVERERERERVVVVVVVV3d3dmZmZVVVVVVVVVVVUzMzMzMzNERERVVVVERERVVVV3d3dVVVVERERVVVVVVVVEREQzMzNERERERERVVVVVVVVVVVVERERVVVVERERVVVVEREREREREREQzMzMzMzNERERVVVVmZmZVVVVERERVVVVVVVVmZmZEREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzNEREREREQzMzMiIiIzMzMiIiIzMzMzMzNERERVVVVEREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIzMzNERERERERERERVVVVEREQzMzNEREQzMzNERERERERVVVVVVVVVVVVVVVVEREREREQzMzMzMzNEREREREREREQzMzNERERERERVVVVVVVVVVVVVVVVVVVVEREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzNERERERERERERERERERERVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVERERERERERERERERVVVVVVVVVVVVVVVVEREREREREREREREREREQzMzMzMzMzMzMzMzNEREQzMzNERERERERERERERERERERVVVVmZmZVVVVVVVVEREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVEREQzMzMzMzMzMzMzMzNERERVVVV3d3dmZmZEREQzMzMzMzMzMzMiIiJERESIiIiIiIhmZmZmZmZmZmZmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZ3d3dmZmZEREQiIiIzMzNVVVWIiIh3d3d3d3d3d3dmZmZ3d3dmZmZEREREREREREQzMzNEREQzMzMzMzMiIiIiIiIzMzNVVVVmZmZ3d3d3d3eIiIiIiIh3d3d3d3dmZmZmZmZVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVEREQzMzNEREQzMzMzMzMzMzMzMzNEREQzMzNEREREREQzMzNEREQzMzMzMzNERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVEREREREQzMzMzMzNERERERERERERVVVVVVVVmZmZVVVVERERVVVVmZmZmZmZVVVV3d3eIiIiZmZmZmZmIiIh3d3eIiIjMzMzMzMyqqqpVVVUiIiJERESqqqqqqqp3d3dVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERmZmZVVVVVVVVVVVVVVVVmZmZVVVVERERVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZ3d3dmZmZVVVV3d3d3d3eIiIh3d3dmZmZVVVVERERVVVVERERVVVVVVVVmZmZmZmZmZmZmZmZ3d3dmZmZmZmZ3d3eZmZmIiIiIiIiIiIiIiIh3d3dmZmZ3d3eIiIh3d3eIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3eIiIiZmZmZmZl3d3dmZmZmZmZmZmZ3d3d3d3dmZmZmZmZmZmZERERERERmZmZ3d3eqqqq7u7uZmZl3d3dVVVVVVVVEREQzMzNEREREREQzMzNERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZ3d3dmZmZmZmZmZmaIiIiqqqqZmZmZmZm7u7vd3d3MzMyIiIhmZmZmZmZVVVVVVVVmZmZ3d3dmZmZmZmZVVVVVVVVVVVV3d3eIiIjMzMy7u7vMzMy7u7uqqqqIiIiIiIiIiIiIiIiIiIh3d3d3d3dVVVVVVVVEREREREQzMzMzMzMiIiIzMzMzMzMzMzNEREQzMzMzMzMzMzNEREREREQzMzNERERVVVVVVVVmZmZ3d3eZmZm7u7vu7u7///////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////7u7u7u7u7u7u7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMu7u7u7u7u7u7qqqqmZmZiIiImZmZd3d3d3d3iIiImZmZmZmZiIiId3d3iIiIiIiIiIiImZmZmZmZmZmZd3d3mZmZmZmZiIiIiIiIiIiIiIiId3d3iIiIiIiId3d3d3d3iIiId3d3d3d3ZmZmd3d3ZmZmZmZmZmZmVVVVZmZmZmZmVVVVVVVVZmZmVVVVZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVREREREREVVVVVVVVREREREREVVVVREREREREREREREREREREREREREREMzMzREREMzMzREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzVVVVREREREREREREREREREREREREREREREREREREREREREREVVVVVVVVREREREREREREREREREREVVVVZmZmd3d3ZmZmVVVVVVVVVVVVd3d3iIiIiIiIiIiIiIiIZmZmVVVVZmZmd3d3ZmZmZmZmiIiId3d3ZmZmiIiIiIiIiIiId3d3d3d3iIiImZmZd3d3VVVVVVVVd3d3d3d3VVVVVVVVVVVVd3d3ZmZmVVVVVVVVVVVVREREREREREREZmZmmZmZiIiIqqqqzMzMzMzMu7u7qqqqu7u7qqqqu7u7mZmZmZmZmZmZiIiId3d3iIiIiIiImZmZmZmZd3d3mZmZu7u7zMzMu7u7mZmZiIiIiIiIiIiId3d3d3d3d3d3d3d3iIiImZmZmZmZiIiIZmZmVVVVREREREREMzMzZmZmqqqqu7u7qqqqqqqqqqqqmZmZiIiIiIiIiIiIiIiId3d3d3d3mZmZiIiIiIiId3d3VVVVREREVVVVZmZmqqqqu7u7u7u7u7u7qqqqqqqqzMzMzMzMu7u7u7u7u7u7u7u7u7u7qqqqiIiId3d3VVVVREREVVVVd3d3mZmZmZmZmZmZmZmZmZmZmZmZzMzMu7u7qqqqqqqqmZmZmZmZd3d3ZmZmZmZmREREVVVVd3d3iIiIiIiId3d3ZmZmZmZmZmZmd3d3mZmZiIiIiIiIiIiId3d3d3d3iIiIZmZmVVVVREREVVVVd3d3d3d3iIiId3d3d3d3d3d3iIiIiIiIqqqqiIiIZmZmd3d3d3d3iIiId3d3VVVVMzMzVVVVd3d3iIiIiIiId3d3iIiIiIiIqqqqmZmZmZmZmZmZmZmZd3d3ZmZmZmZmVVVVd3d3qqqqmZmZmZmZmZmZiIiIiIiIiIiIiIiImZmZiIiIiIiIiIiId3d3d3d3ZmZmVVVVZmZmd3d3iIiImZmZmZmZmZmZmZmZmZmZmZmZmZmZiIiIiIiIu7u7u7u7qqqqqqqqu7u7qqqqiIiId3d3ZmZmZmZmZmZmd3d3d3d3iIiIiIiId3d3ZmZmd3d3iIiImZmZmZmZd3d3ZmZmVVVVVVVVVVVVd3d3ZmZmVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVd3d3iIiIiIiId3d3iIiIqqqqqqqqd3d3ZmZmVVVVREREVVVVVVVVZmZmZmZmiIiImZmZiIiIqqqqqqqqd3d3iIiIiIiIiIiIZmZmiIiImZmZmZmZmZmZd3d3d3d3ZmZmZmZmZmZmZmZmd3d3d3d3iIiIiIiImZmZmZmZiIiIiIiIZmZmZmZmZmZmiIiId3d3d3d3ZmZmd3d3ZmZmREREREREREREREREREREVVVVVVVVVVVVVVVVREREVVVVREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzREREZmZmZmZmVVVVREREREREREREVVVVREREREREd3d3iIiIZmZmZmZmd3d3d3d3ZmZmREREREREREREVVVVZmZmVVVVVVVVVVVVVVVVREREMzMzREREMzMzVVVVZmZmVVVVREREREREREREVVVVREREMzMzREREREREVVVVREREVVVVREREREREREREREREREREREREREREMzMzREREREREZmZmZmZmVVVVVVVVREREREREVVVVREREREREMzMzREREREREMzMzMzMzMzMzREREMzMzMzMzIiIiMzMzIiIiMzMzIiIiMzMzVVVVVVVVREREREREMzMzMzMzMzMzIiIiIiIiMzMzREREIiIiMzMzIiIiMzMzREREREREREREIiIiMzMzIiIiMzMzIiIiMzMzREREREREREREVVVVVVVVVVVVREREREREMzMzREREMzMzREREREREVVVVREREREREREREIiIiMzMzREREREREMzMzMzMzMzMzREREVVVVVVVVREREVVVVREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzIiIiMzMzMzMzIiIiIiIiIiIiMzMzREREREREREREREREREREREREVVVVREREREREMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREREREREREREREREREVVVVVVVVVVVVREREVVVVREREREREREREREREMzMzREREREREREREMzMzMzMzREREREREREREREREREREREREVVVVZmZmVVVVVVVVVVVVREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzMzMzIiIiMzMzREREREREVVVVVVVVMzMzMzMzREREMzMzMzMzMzMzd3d3d3d3VVVVd3d3d3d3ZmZmVVVVVVVVREREREREVVVVVVVVVVVVZmZmZmZmd3d3ZmZmVVVVMzMzMzMzREREZmZmZmZmVVVVd3d3ZmZmZmZmZmZmREREREREREREREREMzMzREREREREREREMzMzREREREREZmZmd3d3iIiIiIiIiIiId3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVZmZmREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVZmZmVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmVVVVREREREREMzMzREREREREREREMzMzVVVVVVVVVVVVZmZmREREVVVVZmZmZmZmVVVVZmZmmZmZmZmZmZmZiIiIiIiIZmZmiIiIzMzMzMzMmZmZVVVVMzMzMzMzmZmZqqqqd3d3ZmZmVVVVVVVVVVVVREREVVVVZmZmVVVVVVVVZmZmZmZmREREREREREREREREVVVVZmZmREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3ZmZmd3d3d3d3iIiIqqqqu7u7iIiIZmZmVVVVREREREREVVVVVVVVZmZmVVVVVVVVZmZmVVVVZmZmZmZmZmZmiIiImZmZmZmZmZmZmZmZiIiIiIiIiIiId3d3d3d3iIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3iIiIiIiIZmZmZmZmVVVVVVVVZmZmVVVVZmZmVVVVREREMzMzVVVVd3d3ZmZmZmZmd3d3d3d3ZmZmZmZmVVVVREREVVVVREREREREREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmd3d3iIiIu7u7zMzMzMzMu7u7iIiIVVVVZmZmd3d3VVVVZmZmZmZmd3d3ZmZmVVVVVVVVZmZmZmZmiIiIu7u7qqqqu7u7qqqqmZmZiIiIiIiIiIiImZmZiIiIZmZmZmZmd3d3VVVVREREREREMzMzIiIiIiIiMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREMzMzREREVVVVZmZmZmZmd3d3u7u73d3d7u7u////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7t3d3e7u7u7u7u7u7t3d3e7u7u7u7u7u7t3d3e7u7t3d3e7u7u7u7u7u7t3d3e7u7t3d3d3d3czMzN3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzLu7u8zMzMzMzN3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3e7u7t3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3czMzMzMzLu7u7u7u6qqqqqqqpmZmYiIiJmZmYiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZnd3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVURERFVVVVVVVVVVVURERFVVVURERERERERERERERFVVVURERERERERERERERDMzM0RERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzM0RERERERERERFVVVVVVVWZmZlVVVVVVVURERERERFVVVURERFVVVVVVVVVVVVVVVURERFVVVWZmZlVVVWZmZmZmZnd3d2ZmZmZmZmZmZmZmZnd3d5mZmZmZmZmZmYiIiIiIiHd3d2ZmZnd3d3d3d4iIiKqqqpmZmYiIiIiIiIiIiJmZmYiIiIiIiJmZmaqqqoiIiGZmZlVVVWZmZmZmZmZmZlVVVVVVVWZmZmZmZlVVVURERFVVVURERERERDMzM0RERFVVVXd3d6qqqszMzMzMzLu7u6qqqqqqqqqqqpmZmZmZmZmZmZmZmYiIiHd3d3d3d3d3d3d3d3d3d3d3d4iIiJmZmZmZmbu7u5mZmXd3d4iIiIiIiHd3d2ZmZmZmZnd3d4iIiIiIiIiIiHd3d2ZmZlVVVURERDMzMzMzM2ZmZpmZmaqqqpmZmYiIiJmZmYiIiIiIiIiIiJmZmYiIiIiIiJmZmaqqqpmZmZmZmYiIiFVVVVVVVVVVVWZmZqqqqru7u6qqqpmZmZmZmZmZmaqqqqqqqru7u6qqqqqqqqqqqpmZmYiIiHd3d4iIiFVVVVVVVWZmZnd3d3d3d3d3d4iIiHd3d3d3d4iIiJmZmYiIiGZmZnd3d4iIiHd3d3d3d1VVVWZmZlVVVWZmZnd3d3d3d3d3d4iIiHd3d3d3d4iIiKqqqoiIiIiIiGZmZmZmZmZmZmZmZmZmZmZmZlVVVURERHd3d4iIiJmZmZmZmYiIiHd3d4iIiIiIiIiIiKqqqpmZmXd3d2ZmZmZmZmZmZlVVVURERERERGZmZpmZmZmZmZmZmaqqqoiIiIiIiJmZmYiIiIiIiIiIiIiIiHd3d2ZmZmZmZlVVVXd3d5mZmYiIiHd3d4iIiHd3d3d3d4iIiJmZmYiIiJmZmXd3d3d3d3d3d3d3d2ZmZlVVVVVVVWZmZoiIiIiIiJmZmZmZmYiIiJmZmZmZmZmZmYiIiIiIiJmZmZmZmaqqqqqqqqqqqmZmZlVVVVVVVWZmZmZmZmZmZmZmZnd3d4iIiHd3d3d3d2ZmZlVVVWZmZnd3d4iIiIiIiFVVVVVVVWZmZmZmZoiIiHd3d1VVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVXd3d5mZmZmZmYiIiIiIiJmZmaqqqoiIiGZmZlVVVVVVVVVVVWZmZlVVVXd3d4iIiJmZmZmZmbu7u6qqqpmZmZmZmYiIiHd3d3d3d3d3d5mZmZmZmYiIiHd3d4iIiIiIiHd3d2ZmZmZmZnd3d4iIiJmZmaqqqoiIiIiIiIiIiHd3d1VVVVVVVXd3d2ZmZlVVVWZmZmZmZnd3d2ZmZlVVVURERERERERERDMzM0RERERERFVVVURERFVVVVVVVTMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERERERFVVVWZmZlVVVVVVVWZmZmZmZkRERFVVVXd3d3d3d3d3d3d3d2ZmZmZmZlVVVVVVVVVVVURERFVVVVVVVVVVVTMzM1VVVVVVVURERERERDMzM0RERGZmZnd3d1VVVURERERERERERERERERERERERERERFVVVVVVVURERERERERERERERDMzM0RERERERFVVVURERERERDMzM1VVVWZmZlVVVURERFVVVURERERERERERERERERERDMzM0RERDMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIkRERGZmZkRERERERERERDMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzMyIiIiIiIjMzM0RERFVVVURERERERFVVVWZmZkRERFVVVURERDMzM0RERERERDMzM0RERERERERERERERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERFVVVURERERERERERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzM0RERERERERERFVVVURERERERERERERERERERDMzMzMzMzMzMzMzM0RERDMzMzMzM0RERDMzM0RERERERERERERERERERGZmZlVVVVVVVVVVVURERERERERERERERDMzM0RERDMzM0RERERERDMzMzMzM0RERFVVVURERERERERERFVVVWZmZmZmZlVVVVVVVURERERERERERERERDMzMzMzMzMzM0RERDMzMzMzM0RERFVVVTMzMzMzMzMzM0RERFVVVURERERERDMzM0RERERERDMzM0RERCIiIjMzM2ZmZmZmZlVVVWZmZmZmZkRERERERERERERERERERFVVVVVVVWZmZmZmZnd3d2ZmZnd3d2ZmZkRERCIiIjMzMzMzM1VVVWZmZmZmZnd3d3d3d2ZmZlVVVURERERERERERERERERERERERERERERERERERGZmZmZmZnd3d4iIiJmZmXd3d2ZmZkRERFVVVVVVVVVVVVVVVURERFVVVVVVVVVVVWZmZlVVVVVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERDMzMzMzMyIiIjMzMyIiIjMzMzMzM1VVVWZmZlVVVVVVVURERERERERERFVVVVVVVWZmZkRERDMzMzMzMzMzMzMzM1VVVURERERERERERERERGZmZlVVVVVVVVVVVVVVVVVVVWZmZoiIiJmZmZmZmZmZmYiIiGZmZnd3d3d3d5mZmbu7u5mZmVVVVTMzM0RERJmZmZmZmWZmZlVVVVVVVVVVVURERERERERERFVVVWZmZmZmZnd3d2ZmZkRERERERERERERERFVVVVVVVVVVVVVVVVVVVURERERERGZmZnd3d1VVVXd3d2ZmZnd3d3d3d5mZmYiIiKqqqszMzJmZmXd3d0RERERERERERFVVVVVVVURERFVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVWZmZmZmZnd3d3d3d3d3d3d3d2ZmZnd3d2ZmZmZmZnd3d2ZmZmZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZnd3d1VVVURERFVVVVVVVWZmZlVVVTMzMzMzM0RERERERERERERERFVVVVVVVURERGZmZlVVVVVVVVVVVURERFVVVVVVVWZmZmZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZqqqqszMzN3d3d3d3czMzIiIiFVVVWZmZnd3d2ZmZlVVVWZmZnd3d2ZmZlVVVWZmZnd3d2ZmZmZmZoiIiIiIiJmZmaqqqqqqqoiIiGZmZmZmZpmZmaqqqnd3d2ZmZmZmZlVVVURERDMzMyIiIiIiIjMzMzMzMzMzMzMzM0RERDMzM0RERDMzMzMzMzMzMzMzM0RERFVVVWZmZnd3d6qqqszMzN3d3f///////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3d3d3u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3d3d3d3d3d3d3u7u7d3d3u7u7d3d3d3d3u7u7d3d3d3d3d3d3d3d3d3d3MzMzd3d3MzMzMzMzMzMzMzMy7u7u7u7uqqqqqqqqZmZmZmZmIiIiIiIiIiIiIiIh3d3d3d3dmZmZmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVEREQzMzNERERVVVVERERVVVVERERVVVVERERERERVVVVEREREREQzMzNEREREREREREQzMzNEREREREREREREREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzNEREQzMzMzMzNERERVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZ3d3dmZmZVVVVVVVV3d3d3d3d3d3dmZmZ3d3d3d3dmZmZ3d3eIiIh3d3d3d3eIiIiZmZmqqqqZmZmZmZl3d3d3d3d3d3dmZmZ3d3eZmZmqqqqZmZl3d3eIiIiZmZmZmZmZmZmqqqq7u7uqqqqIiIhmZmZmZmaIiIhmZmZmZmZVVVVmZmZmZmZVVVVVVVVmZmZVVVUzMzNERERERERmZmZmZmaqqqrMzMzMzMy7u7uqqqqZmZmZmZmZmZmIiIiqqqqZmZmZmZmIiIh3d3d3d3dmZmZVVVV3d3eqqqqZmZl3d3eIiIiIiIh3d3eZmZmZmZl3d3dmZmZVVVVmZmaIiIiZmZmZmZl3d3d3d3dmZmZVVVVEREQzMzNmZmaqqqq7u7uIiIiIiIiIiIiIiIiIiIiqqqqqqqqZmZmqqqqqqqqqqqqZmZl3d3d3d3dmZmZERERERERmZmaqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqq7u7uqqqqZmZmIiIh3d3d3d3d3d3dmZmZ3d3d3d3eIiIiIiIiIiIiZmZmZmZmIiIiIiIiIiIh3d3dmZmZ3d3eZmZmZmZmIiIhmZmZVVVVmZmZmZmaIiIiIiIiZmZmIiIiZmZmIiIiZmZmqqqqqqqqIiIiIiIh3d3d3d3d3d3dmZmZmZmZVVVVmZmaIiIiIiIiIiIiZmZmIiIiIiIiZmZmZmZmZmZmZmZmZmZl3d3dmZmZERERVVVVEREQzMzNVVVV3d3eqqqqqqqqqqqqqqqqZmZmIiIiIiIiIiIiZmZl3d3d3d3d3d3dmZmZ3d3dVVVVmZmaIiIiIiIh3d3eIiIiIiIh3d3eIiIiZmZmZmZmIiIh3d3d3d3d3d3d3d3dmZmZVVVVVVVV3d3eIiIiZmZmZmZmIiIiIiIiIiIiZmZmIiIiIiIh3d3d3d3d3d3eZmZmZmZl3d3dmZmZmZmZ3d3dmZmZ3d3dmZmZVVVVVVVVmZmZ3d3d3d3dmZmZVVVVVVVVVVVV3d3dmZmZVVVVmZmZmZmZ3d3d3d3d3d3dVVVVVVVVERERVVVVERERVVVVmZmZmZmZVVVVVVVVERERmZmZ3d3eZmZmqqqqZmZl3d3d3d3eIiIiZmZmZmZl3d3dmZmZVVVVVVVVVVVVVVVV3d3eIiIiIiIiqqqrMzMyqqqqqqqqIiIh3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIh3d3dmZmZmZmaIiIiZmZmIiIiqqqqIiIiIiIiIiIh3d3dVVVVVVVV3d3dmZmZVVVVVVVVVVVVmZmZEREREREREREQzMzMzMzMzMzNERERERERVVVVVVVVEREREREQzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzNVVVVVVVVVVVVmZmZmZmZVVVVERERERERVVVV3d3d3d3d3d3d3d3dmZmZmZmZmZmZVVVVVVVVERERERERVVVVVVVVERERERERERERERERERERERERmZmZ3d3dmZmZEREREREREREREREREREQzMzNEREREREREREREREREREREREREREREREREREQzMzNERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZVVVUzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNVVVVVVVVEREREREQzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzNEREREREQzMzMzMzMzMzNERERmZmZERERERERERERVVVVVVVVERERERERVVVUzMzNEREREREREREQzMzMzMzNEREQzMzNEREQzMzNEREREREQzMzMzMzMzMzMzMzNERERVVVVERERERERVVVVERERERERERERVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMiIiIREREiIiIzMzNEREREREREREREREREREREREREREQzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzNEREQzMzMzMzNERERVVVVVVVVVVVVVVVVVVVVEREREREREREREREQzMzNEREREREQzMzNERERERERERERERERERERERERERERVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVEREREREREREREREQzMzMzMzMzMzMzMzNEREREREREREQzMzNERERVVVVERERVVVVVVVVEREQzMzNEREQzMzNEREQzMzMiIiJ3d3eIiIhVVVVERERERERVVVVVVVVVVVVERERERERERERVVVVVVVVmZmZmZmZmZmZ3d3dmZmZEREQzMzMzMzNERERVVVVmZmZmZmZ3d3d3d3dmZmZVVVVEREREREREREREREQzMzMzMzMzMzNERERVVVVmZmZ3d3d3d3d3d3d3d3d3d3dVVVVERERERERVVVVVVVVERERERERERERVVVVERERVVVVmZmZVVVVEREREREQzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVVVVVVVVVERERERERVVVVERERVVVVmZmZVVVVEREQzMzMzMzMzMzMzMzNERERVVVVVVVVERERERERVVVVERERVVVVVVVVmZmZmZmZ3d3d3d3eIiIiZmZmZmZl3d3dmZmZmZmaIiIiqqqq7u7uZmZlVVVUzMzMzMzOZmZmZmZlmZmZmZmZVVVVERERERERERERVVVVERERVVVVVVVVmZmZVVVVERERVVVVERERVVVVVVVVVVVVVVVVERERVVVVERERERERmZmaIiIh3d3d3d3d3d3dmZmZ3d3eIiIiZmZmZmZmZmZmIiIhmZmZERERVVVVERERVVVVERERERERVVVVVVVVERERVVVVmZmZVVVVERERERERVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVV3d3dmZmZVVVVERERERERERERVVVVmZmZVVVVERERERERERERERERmZmZVVVVERERVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZmZmZ3d3dmZmZ3d3d3d3d3d3dmZmZ3d3eqqqrMzMzd3d3d3d3d3d27u7uIiIh3d3dmZmZVVVVmZmZmZmZ3d3eIiIh3d3d3d3dmZmZVVVV3d3dmZmZ3d3eZmZnMzMy7u7uZmZlmZmZ3d3eZmZmqqqqqqqqIiIhmZmZEREQzMzMzMzMiIiIzMzMzMzMzMzNEREQzMzMzMzNEREREREREREQzMzNERERERERVVVVmZmZ3d3eZmZm7u7vd3d3////////////////u7u7///////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u3d3d7u7u3d3d3d3d7u7u7u7u7u7u3d3d7u7u7u7u7u7u3d3d7u7u7u7u7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7qqqqqqqqqqqqqqqqmZmZmZmZiIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3iIiIiIiIZmZmZmZmVVVVREREMzMzMzMzREREREREREREREREVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREVVVVREREREREVVVVZmZmZmZmZmZmd3d3ZmZmZmZmZmZmmZmZmZmZiIiIiIiId3d3iIiId3d3iIiIqqqqmZmZd3d3iIiImZmZqqqqqqqqmZmZqqqqmZmZiIiIiIiId3d3iIiImZmZmZmZiIiImZmZqqqqmZmZqqqqqqqqqqqqmZmZqqqqd3d3d3d3iIiIZmZmZmZmVVVVZmZmd3d3ZmZmd3d3ZmZmVVVVREREMzMzREREZmZmiIiIu7u7zMzMzMzMu7u7u7u7mZmZiIiId3d3iIiIiIiImZmZmZmZiIiId3d3ZmZmVVVVVVVViIiIqqqqmZmZd3d3d3d3iIiId3d3mZmZmZmZd3d3ZmZmZmZmd3d3d3d3iIiImZmZZmZmVVVVVVVVREREREREMzMzZmZmiIiImZmZmZmZiIiImZmZmZmZmZmZqqqqmZmZmZmZqqqqmZmZiIiId3d3ZmZmREREREREREREREREd3d3u7u73d3dzMzMu7u7qqqqu7u7u7u7mZmZqqqqu7u7qqqqqqqqmZmZiIiId3d3ZmZmd3d3mZmZqqqqqqqqqqqqqqqqqqqqqqqqu7u7qqqqmZmZmZmZd3d3iIiImZmZmZmZd3d3VVVVZmZmd3d3d3d3iIiImZmZmZmZmZmZmZmZmZmZiIiImZmZmZmZmZmZmZmZiIiImZmZd3d3ZmZmZmZmVVVVd3d3iIiId3d3iIiImZmZqqqqqqqqqqqqqqqqmZmZmZmZiIiIVVVVVVVVREREVVVVREREMzMzREREd3d3qqqqu7u7qqqqqqqqmZmZiIiImZmZmZmZiIiId3d3d3d3ZmZmiIiId3d3VVVVZmZmmZmZd3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3iIiId3d3VVVVVVVVVVVVZmZmmZmZqqqqiIiId3d3iIiId3d3iIiIiIiIiIiId3d3d3d3d3d3mZmZmZmZiIiIZmZmZmZmd3d3d3d3d3d3ZmZmZmZmVVVVVVVVZmZmd3d3d3d3VVVVVVVVVVVVd3d3ZmZmZmZmd3d3ZmZmd3d3d3d3ZmZmVVVVZmZmVVVVREREREREVVVVVVVVZmZmZmZmZmZmVVVVd3d3mZmZqqqqqqqqiIiIZmZmiIiIiIiIiIiIqqqqmZmZZmZmZmZmVVVVREREVVVVd3d3d3d3iIiIqqqqu7u7mZmZmZmZiIiId3d3ZmZmZmZmd3d3d3d3mZmZd3d3iIiIiIiIiIiId3d3ZmZmZmZmiIiIiIiImZmZiIiIiIiIiIiIZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREMzMzMzMzREREREREREREREREVVVVREREREREMzMzMzMzMzMzMzMzREREREREMzMzMzMzREREREREVVVVVVVVZmZmVVVVREREREREZmZmiIiId3d3d3d3d3d3ZmZmZmZmd3d3ZmZmVVVVVVVVREREREREVVVVREREREREMzMzREREREREZmZmd3d3d3d3REREREREREREREREREREREREREREREREREREREREREREREREREREZmZmREREREREREREMzMzREREREREREREREREZmZmVVVVVVVVVVVVVVVVVVVVREREREREMzMzREREVVVVMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREZmZmREREREREREREMzMzREREREREMzMzMzMzIiIiMzMzMzMzMzMzREREREREMzMzREREREREMzMzREREMzMzMzMzMzMzREREZmZmREREREREREREVVVVVVVVREREVVVVREREMzMzMzMzVVVVREREMzMzMzMzMzMzMzMzREREREREMzMzMzMzMzMzMzMzIiIiMzMzVVVVVVVVREREREREREREREREVVVVREREREREREREREREMzMzMzMzIiIiMzMzIiIiMzMzREREMzMzMzMzREREMzMzMzMzIiIiIiIiMzMzMzMzREREREREVVVVREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREMzMzMzMzMzMzMzMzMzMzREREVVVVZmZmVVVVVVVVREREREREREREREREREREREREREREREREREREMzMzREREMzMzREREMzMzREREMzMzREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREMzMzREREMzMzMzMzMzMzMzMzMzMzREREREREMzMzREREREREVVVVVVVVVVVVVVVVREREREREMzMzMzMzMzMzMzMzIiIiZmZmd3d3VVVVMzMzREREZmZmZmZmVVVVREREREREREREVVVVVVVVVVVVZmZmZmZmd3d3d3d3REREREREREREREREVVVVZmZmZmZmd3d3iIiId3d3ZmZmREREREREREREREREMzMzMzMzREREREREREREVVVVd3d3d3d3iIiId3d3ZmZmREREREREREREVVVVVVVVREREREREVVVVREREVVVVZmZmZmZmVVVVREREREREMzMzMzMzMzMzIiIiERERIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzVVVVVVVVVVVVREREREREREREREREVVVVREREVVVVVVVVVVVVREREREREMzMzMzMzREREREREREREREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3ZmZmZmZmd3d3iIiId3d3d3d3d3d3mZmZu7u7zMzMmZmZVVVVMzMzREREmZmZmZmZZmZmVVVVREREREREMzMzREREREREVVVVREREREREVVVVZmZmREREREREREREREREVVVVREREREREREREREREREREREREZmZmiIiIiIiIiIiImZmZd3d3VVVViIiIiIiId3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVREREVVVVVVVVVVVVVVVVREREREREREREVVVVREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVd3d3ZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVREREREREREREREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVZmZmZmZmVVVVZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmd3d3qqqqzMzM3d3d3d3d3d3d3d3du7u7d3d3ZmZmVVVVVVVVZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmd3d3iIiIu7u73d3du7u7mZmZiIiIiIiImZmZmZmZqqqqiIiIVVVVREREMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzMzMzREREREREVVVVZmZmmZmZzMzM3d3d////////////////////////////////////7u7u////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////+7u7t3d3e7u7u7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3czMzMzMzLu7u7u7u7u7u6qqqqqqqru7u7u7u8zMzLu7u7u7u7u7u7u7u8zMzLu7u7u7u7u7u6qqqqqqqpmZmZmZmYiIiHd3d3d3d2ZmZnd3d2ZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZnd3d3d3d2ZmZkRERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIhERESIiIhERESIiIhERESIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMzMzMyIiIiIiIjMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVVVVVWZmZmZmZmZmZnd3d4iIiIiIiHd3d4iIiJmZmYiIiIiIiJmZmaqqqqqqqoiIiJmZmbu7u7u7u6qqqqqqqqqqqru7u7u7u5mZmYiIiIiIiIiIiJmZmZmZmZmZmaqqqqqqqqqqqqqqqpmZmYiIiIiIiJmZmYiIiIiIiHd3d3d3d2ZmZnd3d2ZmZnd3d3d3d2ZmZlVVVVVVVURERERERFVVVXd3d7u7u93d3czMzMzMzLu7u6qqqoiIiIiIiJmZmZmZmaqqqqqqqpmZmZmZmYiIiHd3d1VVVXd3d4iIiJmZmXd3d3d3d3d3d3d3d4iIiIiIiIiIiJmZmXd3d3d3d3d3d3d3d2ZmZlVVVURERERERERERFVVVURERGZmZpmZmaqqqqqqqqqqqqqqqqqqqpmZmZmZmYiIiKqqqpmZmZmZmaqqqoiIiGZmZmZmZmZmZmZmZlVVVZmZmd3d3czMzLu7u7u7u7u7u6qqqpmZmYiIiLu7u7u7u6qqqpmZmZmZmZmZmXd3d2ZmZoiIiHd3d4iIiLu7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqqqqqqqqqpmZmZmZmYiIiHd3d2ZmZnd3d4iIiHd3d4iIiLu7u6qqqqqqqqqqqpmZmZmZmZmZmZmZmaqqqoiIiHd3d4iIiHd3d3d3d3d3d1VVVVVVVXd3d3d3d4iIiKqqqpmZmZmZmZmZmYiIiIiIiIiIiHd3d1VVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d6qqqqqqqnd3d5mZmYiIiIiIiIiIiHd3d3d3d2ZmZnd3d3d3d5mZmWZmZlVVVXd3d5mZmXd3d2ZmZnd3d4iIiIiIiIiIiIiIiIiIiHd3d3d3d5mZmXd3d3d3d1VVVWZmZnd3d3d3d4iIiKqqqoiIiIiIiHd3d4iIiHd3d4iIiIiIiIiIiIiIiHd3d5mZmZmZmYiIiIiIiHd3d4iIiIiIiGZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZnd3d4iIiHd3d3d3d2ZmZmZmZmZmZnd3d3d3d2ZmZmZmZlVVVURERERERERERFVVVVVVVVVVVVVVVVVVVYiIiKqqqqqqqoiIiHd3d2ZmZnd3d4iIiIiIiJmZmZmZmXd3d3d3d2ZmZlVVVVVVVVVVVXd3d5mZmaqqqpmZmYiIiIiIiHd3d3d3d1VVVVVVVXd3d4iIiIiIiHd3d3d3d3d3d4iIiHd3d1VVVWZmZnd3d4iIiJmZmYiIiIiIiIiIiHd3d1VVVURERGZmZmZmZlVVVVVVVWZmZlVVVXd3d2ZmZnd3d2ZmZkRERDMzM0RERERERERERDMzM0RERFVVVVVVVURERERERDMzM0RERDMzM0RERDMzMzMzM0RERDMzM0RERERERFVVVVVVVVVVVVVVVWZmZoiIiIiIiHd3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVURERERERERERFVVVURERERERDMzMzMzMzMzM0RERIiIiGZmZlVVVURERERERFVVVURERERERERERERERERERERERERERFVVVURERFVVVURERERERDMzMzMzMzMzMzMzMzMzM1VVVWZmZlVVVVVVVVVVVWZmZlVVVURERERERDMzM0RERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVWZmZlVVVURERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzM0RERDMzMyIiIkRERERERERERERERFVVVVVVVURERDMzM1VVVWZmZjMzM1VVVVVVVURERDMzM0RERERERDMzM0RERDMzMzMzMzMzMzMzMzMzM0RERFVVVTMzMzMzMzMzM0RERFVVVURERERERERERERERERERERERERERFVVVURERERERDMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzMzMzMzMzMzMzM0RERCIiIjMzM1VVVURERERERFVVVURERERERERERERERERERDMzMzMzM0RERDMzMzMzMzMzM0RERERERERERDMzM0RERDMzMzMzMzMzMzMzM1VVVWZmZlVVVVVVVURERERERERERERERERERFVVVURERERERERERERERDMzM0RERERERERERDMzMzMzMzMzM0RERFVVVURERERERFVVVVVVVURERDMzM0RERERERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERDMzMzMzM0RERFVVVXd3d4iIiHd3d0RERERERDMzMyIiIiIiIkRERGZmZlVVVURERERERGZmZmZmZlVVVURERERERERERERERERERFVVVVVVVXd3d4iIiHd3d1VVVURERERERDMzM0RERGZmZmZmZnd3d5mZmYiIiHd3d1VVVURERERERERERERERDMzM2ZmZkRERDMzM0RERGZmZmZmZmZmZoiIiGZmZmZmZlVVVURERFVVVURERFVVVURERERERFVVVVVVVVVVVWZmZmZmZkRERERERDMzMzMzMyIiIhERESIiIhERERERESIiIiIiIiIiIjMzMzMzM0RERDMzMyIiIjMzMzMzMzMzM0RERFVVVVVVVURERERERERERERERERERERERERERFVVVVVVVURERFVVVURERERERERERERERERERFVVVVVVVURERFVVVURERFVVVWZmZnd3d3d3d1VVVVVVVVVVVXd3d3d3d3d3d3d3d3d3d4iIiLu7u6qqqoiIiGZmZjMzMzMzM3d3d3d3d2ZmZlVVVURERERERERERERERERERFVVVURERERERFVVVWZmZkRERDMzM0RERDMzM0RERERERERERERERERERERERERERGZmZoiIiIiIiIiIiKqqqpmZmXd3d2ZmZmZmZlVVVWZmZmZmZnd3d1VVVWZmZoiIiGZmZmZmZmZmZoiIiJmZmYiIiFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERERERFVVVURERERERERERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVURERERERERERFVVVWZmZmZmZnd3d2ZmZlVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVURERFVVVVVVVWZmZmZmZlVVVWZmZmZmZnd3d2ZmZmZmZnd3d3d3d3d3d7u7u93d3d3d3czMzMzMzKqqqoiIiGZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZnd3d2ZmZlVVVWZmZpmZmaqqqru7u5mZmZmZmaqqqqqqqpmZmYiIiHd3d2ZmZlVVVURERDMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVVVVVURERERERDMzM0RERERERERERFVVVXd3d6qqqt3d3e7u7v///////////////////////////////////////////+7u7v///////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3MzMzMzMy7u7u7u7uqqqqZmZmZmZmZmZmZmZmqqqq7u7vMzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3MzMzMzMy7u7vMzMy7u7uqqqqZmZmIiIh3d3d3d3dmZmZmZmZmZmZ3d3d3d3d3d3d3d3eIiIiIiIiZmZmIiIh3d3dmZmZVVVVEREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNEREQzMzMiIiIzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzNERERVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVV3d3dmZmaIiIiZmZmqqqqqqqqqqqqZmZmqqqqqqqqqqqqZmZmqqqq7u7uZmZmIiIiIiIiIiIh3d3eIiIiIiIiIiIiZmZmqqqqqqqqqqqqZmZl3d3d3d3eIiIiZmZmIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3dVVVVERERERERERERERERmZmaqqqrMzMzMzMzMzMzMzMyqqqq7u7uqqqqqqqq7u7u7u7uqqqqZmZmZmZmIiIhVVVVmZmZ3d3eZmZmZmZmIiIiqqqqZmZl3d3d3d3eIiIiIiIh3d3eIiIiIiIh3d3eIiIh3d3dVVVVERERVVVVVVVVVVVVVVVWIiIi7u7uqqqqZmZmZmZmqqqqZmZmIiIiIiIiZmZmZmZmZmZmZmZmqqqqIiIhmZmZ3d3eZmZl3d3dmZmaZmZnd3d3d3d27u7u7u7uqqqqZmZmIiIiqqqq7u7u7u7uqqqqZmZmZmZmIiIh3d3eIiIiIiIhmZmaIiIi7u7vMzMy7u7u7u7vMzMy7u7uqqqq7u7uqqqqqqqqZmZmZmZmZmZl3d3eIiIiZmZl3d3dmZmaZmZnMzMy7u7u7u7uqqqqZmZmZmZmqqqqZmZmqqqqIiIh3d3d3d3d3d3d3d3dmZmZVVVVVVVV3d3eIiIh3d3d3d3eIiIiIiIiIiIh3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3d3d3eIiIiZmZmIiIh3d3eIiIiIiIiIiIh3d3eIiIiIiIiIiIhmZmZVVVV3d3d3d3d3d3d3d3eIiIh3d3d3d3d3d3dmZmZ3d3d3d3d3d3eZmZmZmZmIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhmZmZmZmaIiIiIiIh3d3d3d3dmZmZ3d3eIiIiIiIiIiIiZmZmZmZmZmZmqqqqZmZmIiIh3d3eIiIhmZmZ3d3d3d3dmZmZ3d3dmZmZ3d3d3d3dmZmZVVVV3d3eZmZl3d3dmZmZmZmZmZmZVVVVVVVV3d3d3d3d3d3dmZmZVVVVVVVVEREQzMzNERERERERVVVVVVVV3d3eqqqqqqqqIiIh3d3d3d3dmZmZ3d3eZmZmIiIiIiIh3d3eIiIiIiIhmZmZmZmZVVVVmZmaIiIiZmZmqqqqZmZmqqqqIiIhmZmZ3d3dmZmZmZmZ3d3eZmZmIiIh3d3dmZmZ3d3d3d3dmZmZVVVVmZmZ3d3eIiIiqqqqIiIiIiIiIiIh3d3dmZmZVVVVmZmZ3d3dVVVVVVVVmZmZmZmaIiIiIiIh3d3dVVVVVVVVERERERERERERERERERERERERVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERVVVVVVVVERERVVVV3d3eIiIiIiIh3d3d3d3dmZmZVVVVVVVVVVVVERERERERERERERERVVVVmZmZVVVVEREREREQzMzMzMzNERER3d3dmZmZVVVVVVVVVVVVERERERERVVVVERERERERERERERERVVVVVVVVEREREREREREREREREREQzMzMiIiIzMzNERERmZmZmZmZmZmZ3d3dmZmZ3d3dEREREREQzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzNERERERERVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIzMzMzMzMzMzMzMzNVVVVVVVVVVVVVVVVERERERERVVVVVVVVEREREREREREREREQzMzNEREREREQzMzNEREQzMzNEREQzMzMzMzMzMzMzMzNVVVVEREQzMzMzMzMzMzNVVVVVVVVEREREREREREREREREREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzNEREREREQzMzMzMzNERERVVVVERERERERVVVVEREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNEREREREREREQzMzMzMzMiIiIzMzNVVVVVVVVVVVVERERVVVVERERERERERERERERERERERERERERERERVVVVEREREREQzMzNEREREREQzMzMiIiJERERERERERERVVVVEREREREREREREREREREQzMzNEREQzMzNEREREREREREREREREREREREREREQzMzMzMzMzMzNmZmaIiIiqqqqIiIhVVVVEREQzMzMiIiIiIiJVVVVVVVVVVVVERERVVVVERERmZmZVVVVERERERERVVVVVVVVVVVVVVVVVVVVmZmaIiIh3d3dVVVVERERERERERERERERmZmZmZmaIiIiZmZmZmZl3d3dVVVVVVVVEREREREQzMzMzMzNERERERERERERVVVVVVVVERERVVVV3d3d3d3d3d3dmZmZVVVVVVVVVVVVVVVVmZmZVVVVERERERERERERVVVVmZmZVVVUzMzMzMzMiIiIiIiIiIiIiIiIiIiIREREREREiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVEREREREQzMzNEREQzMzNERERVVVVERERVVVVVVVVERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVERERVVVVmZmZ3d3dmZmZVVVVERERmZmZ3d3dmZmaIiIh3d3d3d3eIiIiqqqqqqqqIiIhmZmYzMzMzMzNmZmaIiIhmZmZmZmZVVVVERERERERERERVVVVVVVVVVVVERERERERVVVVVVVVERERERERERERVVVVERERERERERERERERERERVVVVVVVVmZmZ3d3eZmZmZmZmZmZmZmZl3d3dVVVVVVVV3d3d3d3dmZmZVVVV3d3eZmZl3d3dVVVVmZmaZmZm7u7uZmZlVVVVmZmZmZmZmZmZ3d3d3d3d3d3dmZmZmZmZVVVVmZmZmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVERERVVVVVVVVVVVVmZmZ3d3eIiIh3d3dVVVVmZmZmZmZVVVVVVVVERERVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZ3d3dmZmZmZmZ3d3d3d3eZmZnMzMzd3d3MzMy7u7uZmZl3d3dmZmZmZmZmZmZ3d3dmZmZVVVVmZmZ3d3dmZmZmZmZVVVVmZmZ3d3eIiIiZmZmZmZmZmZnMzMyqqqp3d3dmZmZ3d3d3d3dEREQzMzMzMzMzMzNEREQzMzNERERERER3d3eZmZlmZmZVVVVERERERERERERERERVVVVmZmaqqqrd3d3///////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////3d3d3d3d3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u3d3d3d3d7u7u3d3d3d3d3d3dzMzM3d3d3d3dzMzMzMzMzMzMu7u7qqqqqqqqmZmZmZmZqqqqmZmZqqqqmZmZmZmZu7u7u7u7zMzMzMzM3d3dzMzM3d3dzMzM3d3dzMzM3d3dzMzMzMzMzMzMzMzMu7u7u7u7mZmZiIiId3d3d3d3iIiIiIiIiIiIiIiIiIiImZmZmZmZmZmZmZmZiIiId3d3ZmZmVVVVREREREREREREREREREREREREREREMzMzMzMzREREREREVVVVVVVVREREREREMzMzMzMzREREREREMzMzREREREREMzMzREREREREREREREREMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREREREREREMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREMzMzREREREREREREREREREREMzMzMzMzMzMzREREREREVVVVVVVVZmZmZmZmVVVVVVVVVVVVZmZmVVVVVVVVREREVVVVVVVVZmZmVVVVVVVVZmZmZmZmiIiIiIiImZmZiIiIiIiId3d3iIiImZmZiIiImZmZiIiId3d3d3d3d3d3d3d3d3d3iIiIiIiIZmZmZmZmmZmZqqqqqqqqqqqqd3d3ZmZmd3d3mZmZiIiIiIiId3d3d3d3d3d3d3d3mZmZiIiId3d3d3d3VVVVVVVVREREREREd3d3qqqqzMzMzMzMzMzMzMzMqqqqqqqqqqqqu7u7mZmZqqqqmZmZiIiIiIiIZmZmZmZmd3d3d3d3mZmZzMzMqqqqqqqqmZmZiIiIiIiId3d3iIiIiIiId3d3d3d3d3d3iIiIiIiIVVVVVVVVVVVVVVVVREREVVVVmZmZu7u7qqqqmZmZiIiImZmZiIiId3d3d3d3iIiIiIiIiIiImZmZmZmZiIiIZmZmiIiIqqqqd3d3ZmZmmZmZzMzMzMzMzMzMqqqqqqqqmZmZmZmZqqqqu7u7qqqqu7u7qqqqqqqqmZmZmZmZmZmZmZmZmZmZqqqqqqqqu7u7qqqqu7u7u7u7qqqqu7u7u7u7qqqqqqqqqqqqmZmZmZmZiIiImZmZiIiIiIiIiIiIqqqqu7u7u7u7u7u7mZmZmZmZmZmZmZmZmZmZmZmZiIiId3d3ZmZmd3d3d3d3d3d3ZmZmZmZmd3d3iIiId3d3ZmZmZmZmiIiIiIiIiIiIiIiId3d3ZmZmd3d3d3d3d3d3mZmZmZmZiIiIiIiId3d3d3d3d3d3iIiId3d3d3d3iIiIiIiId3d3d3d3ZmZmZmZmd3d3mZmZiIiIiIiId3d3ZmZmd3d3d3d3d3d3ZmZmd3d3iIiImZmZiIiIiIiIiIiIiIiIiIiImZmZqqqqmZmZZmZmZmZmVVVVZmZmd3d3ZmZmVVVVZmZmZmZmd3d3d3d3mZmZmZmZmZmZmZmZqqqqiIiId3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3ZmZmd3d3mZmZqqqqd3d3VVVVREREVVVVVVVVZmZmd3d3d3d3d3d3ZmZmVVVVVVVVREREMzMzREREREREVVVVZmZmmZmZqqqqmZmZmZmZmZmZd3d3d3d3d3d3qqqqiIiId3d3ZmZmZmZmd3d3iIiIZmZmd3d3d3d3iIiImZmZmZmZqqqqqqqqiIiIZmZmd3d3iIiId3d3d3d3mZmZmZmZZmZmVVVVZmZmZmZmVVVVVVVVZmZmZmZmiIiIqqqqmZmZiIiId3d3d3d3VVVVZmZmZmZmZmZmVVVVVVVVZmZmZmZmd3d3d3d3ZmZmZmZmVVVVVVVVREREREREVVVVREREd3d3ZmZmVVVVREREREREREREREREMzMzMzMzMzMzMzMzREREREREMzMzREREVVVVVVVVMzMzREREd3d3d3d3d3d3d3d3d3d3ZmZmVVVVVVVVVVVVREREVVVVREREREREVVVVVVVVVVVVREREREREREREMzMzVVVVZmZmZmZmVVVVVVVVVVVVREREVVVVREREREREVVVVVVVVREREVVVVVVVVVVVVREREREREREREREREMzMzMzMzIiIiREREZmZmZmZmZmZmZmZmd3d3VVVVREREREREREREREREREREMzMzMzMzREREMzMzMzMzIiIiMzMzMzMzMzMzIiIiMzMzIiIiMzMzREREVVVVVVVVVVVVREREMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzREREREREZmZmZmZmVVVVVVVVREREVVVVREREMzMzREREREREREREREREREREMzMzREREMzMzREREMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREREREREREREREREREREREREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzMzMzREREMzMzREREZmZmVVVVVVVVVVVVREREMzMzREREVVVVREREMzMzREREMzMzREREMzMzREREMzMzMzMzREREREREREREREREMzMzIiIiMzMzMzMzVVVVVVVVREREREREREREREREREREREREREREREREVVVVREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzREREVVVVREREREREVVVVREREMzMzMzMzREREMzMzREREMzMzREREREREREREREREREREVVVVREREZmZmZmZmVVVVd3d3d3d3iIiIZmZmREREMzMzIiIiIiIiZmZmd3d3VVVVREREREREREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVd3d3iIiIiIiId3d3VVVVREREREREREREREREVVVVZmZmiIiIqqqqmZmZd3d3ZmZmVVVVVVVVMzMzREREMzMzMzMzMzMzMzMzREREREREREREREREVVVVd3d3d3d3VVVVREREVVVVVVVVVVVVVVVVVVVVREREREREREREVVVVREREVVVVREREIiIiMzMzMzMzIiIiIiIiIiIiERERIiIiERERIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzVVVVVVVVVVVVREREREREREREMzMzREREREREVVVVREREREREVVVVREREVVVVVVVVREREREREREREREREVVVVVVVVREREVVVVVVVVVVVVZmZmZmZmVVVVVVVVREREVVVVd3d3ZmZmd3d3iIiIiIiId3d3qqqqu7u7mZmZZmZmREREIiIid3d3iIiId3d3VVVVZmZmVVVVREREMzMzREREZmZmVVVVREREREREVVVVZmZmVVVVVVVVREREVVVVREREREREVVVVREREREREREREREREd3d3d3d3iIiIqqqqqqqqmZmZiIiIZmZmVVVVd3d3d3d3ZmZmVVVVd3d3qqqqd3d3ZmZmiIiIqqqqu7u7iIiIZmZmVVVVZmZmZmZmZmZmd3d3mZmZmZmZd3d3ZmZmd3d3d3d3d3d3d3d3ZmZmVVVVZmZmVVVVZmZmd3d3d3d3VVVVZmZmZmZmVVVVZmZmZmZmVVVVVVVVVVVVREREZmZmVVVVZmZmd3d3mZmZqqqqiIiIZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3iIiIqqqqzMzM3d3du7u7qqqqiIiIZmZmZmZmVVVVd3d3ZmZmd3d3ZmZmZmZmZmZmZmZmVVVVVVVVZmZmZmZmiIiImZmZu7u7zMzMmZmZZmZmZmZmiIiImZmZZmZmREREMzMzREREMzMzREREVVVVd3d3d3d3d3d3ZmZmREREREREVVVVVVVVZmZmZmZmiIiIzMzM////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7u7u7u7u7u7u7t3d3d3d3d3d3e7u7u7u7t3d3d3d3d3d3czMzMzMzMzMzLu7u8zMzMzMzN3d3czMzKqqqqqqqqqqqpmZmaqqqqqqqru7u7u7u7u7u7u7u7u7u6qqqru7u6qqqru7u7u7u7u7u8zMzLu7u7u7u8zMzMzMzMzMzMzMzMzMzMzMAP//AADMzMzMu7u7u7u7u7u7qqqqqqqqqqqqqqqqu7u7qqqqmZmZiIiImZmZmZmZiIiIiIiId3d3d3d3iIiId3d3ZmZmZmZmd3d3ZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREREREMzMzREREREREREREREREMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzREREVVVVVVVVREREREREREREREREVVVVREREREREVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmVVVVd3d3d3d3ZmZmVVVVZmZmZmZmZmZmiIiImZmZiIiIiIiId3d3d3d3iIiImZmZiIiId3d3iIiId3d3d3d3iIiIiIiId3d3d3d3ZmZmVVVVVVVVREREVVVVd3d3u7u7zMzMzMzMzMzMzMzMu7u7mZmZqqqqu7u7qqqqmZmZqqqqmZmZd3d3ZmZmd3d3d3d3ZmZmmZmZzMzMqqqqmZmZiIiIiIiIiIiIiIiId3d3d3d3d3d3iIiIiIiId3d3ZmZmVVVVd3d3iIiIVVVVVVVVZmZmmZmZu7u7qqqqmZmZiIiIiIiIiIiIiIiId3d3d3d3iIiId3d3iIiIiIiIiIiId3d3d3d3iIiIiIiId3d3mZmZzMzM3d3du7u7mZmZiIiImZmZqqqqzMzMqqqqqqqqmZmZmZmZmZmZqqqqqqqqu7u7zMzMzMzMu7u7qqqqqqqqmZmZqqqqqqqqu7u7qqqqqqqqqqqqiIiImZmZmZmZmZmZqqqqzMzMu7u7qqqqqqqqqqqqmZmZqqqqmZmZiIiIiIiImZmZmZmZmZmZiIiIiIiId3d3d3d3ZmZmd3d3mZmZmZmZd3d3d3d3iIiIiIiIVVVVVVVVd3d3mZmZiIiIiIiId3d3ZmZmiIiIiIiImZmZmZmZmZmZiIiIiIiId3d3d3d3d3d3d3d3ZmZmiIiIiIiId3d3d3d3d3d3d3d3iIiImZmZmZmZiIiIiIiId3d3ZmZmVVVVZmZmd3d3ZmZmd3d3iIiIiIiIiIiIiIiIqqqqmZmZmZmZqqqqmZmZd3d3ZmZmd3d3iIiId3d3d3d3d3d3ZmZmVVVVZmZmVVVVZmZmmZmZqqqqqqqqqqqqmZmZiIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmd3d3d3d3iIiImZmZd3d3d3d3ZmZmVVVVVVVVVVVVVVVVd3d3d3d3d3d3d3d3ZmZmVVVVREREREREREREREREZmZmmZmZqqqqqqqqmZmZmZmZmZmZd3d3ZmZmd3d3iIiId3d3d3d3ZmZmZmZmZmZmZmZmd3d3iIiId3d3d3d3mZmZmZmZmZmZmZmZiIiId3d3ZmZmd3d3d3d3ZmZmmZmZiIiIZmZmd3d3ZmZmZmZmZmZmVVVVZmZmd3d3mZmZqqqqqqqqd3d3d3d3ZmZmREREZmZmd3d3ZmZmVVVVZmZmd3d3ZmZmVVVVZmZmVVVVREREREREVVVVVVVVVVVVVVVVVVVVZmZmVVVVREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREMzMzREREVVVVVVVVZmZmMzMzREREVVVVd3d3d3d3ZmZmZmZmd3d3ZmZmVVVVREREVVVVVVVVVVVVREREREREREREREREREREREREREREREREVVVVZmZmVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREREREREREMzMzMzMzMzMzVVVVVVVVREREREREVVVVREREREREMzMzMzMzMzMzREREREREVVVVREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiMzMzZmZmVVVVVVVVVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzMzMzREREMzMzMzMzMzMzZmZmVVVVVVVVVVVVVVVVREREREREREREREREREREREREREREREREREREMzMzREREMzMzMzMzREREMzMzMzMzMzMzMzMzREREREREVVVVVVVVVVVVVVVVREREREREVVVVREREREREREREVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzMzMzMzMzMzMzREREVVVVVVVVVVVVREREVVVVVVVVREREMzMzREREREREREREREREMzMzREREREREREREMzMzMzMzMzMzREREMzMzMzMzIiIiIiIiMzMzVVVVREREREREREREVVVVREREVVVVVVVVREREREREREREREREREREREREREREREREMzMzREREREREMzMzREREMzMzREREREREVVVVREREREREREREREREREREMzMzREREREREREREREREVVVVREREREREVVVVZmZmVVVVZmZmd3d3ZmZmZmZmZmZmd3d3d3d3ZmZmMzMzIiIiIiIiZmZmd3d3VVVVREREVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVd3d3iIiId3d3VVVVREREREREREREREREREREVVVVZmZmmZmZqqqqmZmZd3d3ZmZmZmZmREREREREMzMzMzMzMzMzIiIiMzMzMzMzREREREREREREREREVVVVVVVVREREVVVVVVVVVVVVVVVVREREREREREREREREREREREREREREVVVVREREMzMzMzMzMzMzIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzREREREREREREVVVVVVVVVVVVREREMzMzREREREREREREVVVVVVVVREREREREVVVVREREVVVVREREREREREREREREVVVVVVVVREREVVVVREREVVVVZmZmZmZmVVVVVVVVREREREREZmZmd3d3d3d3d3d3iIiIiIiImZmZmZmZqqqqqqqqZmZmMzMzMzMzVVVVmZmZd3d3ZmZmZmZmVVVVMzMzREREREREVVVVVVVVREREREREREREZmZmZmZmZmZmVVVVREREREREVVVVVVVVVVVVREREREREVVVVd3d3d3d3d3d3mZmZmZmZiIiIZmZmZmZmVVVVVVVVVVVVZmZmVVVVZmZmd3d3d3d3iIiImZmZmZmZqqqqd3d3REREVVVVZmZmd3d3d3d3ZmZmiIiIu7u7mZmZZmZmd3d3d3d3iIiIiIiId3d3ZmZmVVVVREREd3d3qqqqd3d3VVVVd3d3ZmZmREREREREZmZmZmZmVVVVVVVVZmZmZmZmVVVVZmZmmZmZmZmZqqqqd3d3VVVVVVVVVVVVVVVVREREVVVVVVVVZmZmZmZmZmZmZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3ZmZmd3d3iIiIiIiIiIiIqqqqiIiImZmZiIiIZmZmVVVVVVVVZmZmZmZmZmZmd3d3d3d3ZmZmVVVVREREVVVVZmZmd3d3mZmZzMzM3d3dqqqqZmZmVVVVZmZmiIiIqqqqZmZmREREREREREREMzMzREREVVVVd3d3d3d3REREREREREREVVVVVVVVVVVVd3d3iIiIzMzM7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////+7u7v///+7u7u7u7u7u7t3d3e7u7t3d3d3d3czMzLu7u7u7u8zMzN3d3d3d3czMzMzMzLu7u7u7u8zMzMzMzMzMzLu7u8zMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u8zMzMzMzMzMzMzMzMzMzN3d3czMzMzMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzLu7u7u7u6qqqpmZmZmZmZmZmYiIiIiIiIiIiJmZmZmZmYiIiIiIiIiIiHd3d3d3d3d3d5mZmYiIiHd3d3d3d3d3d3d3d4iIiIiIiHd3d2ZmZnd3d5mZmYiIiHd3d4iIiJmZmYiIiIiIiJmZmYiIiHd3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d4iIiHd3d4iIiIiIiIiIiHd3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVURERERERERERDMzM0RERDMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMyIiIiIiIjMzMyIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIjMzM0RERERERERERERERERERFVVVURERFVVVWZmZnd3d2ZmZlVVVURERGZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZlVVVVVVVURERGZmZoiIiIiIiIiIiHd3d3d3d5mZmZmZmYiIiJmZmZmZmXd3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVWZmZlVVVURERERERFVVVYiIiKqqqszMzMzMzMzMzN3d3bu7u7u7u7u7u8zMzKqqqpmZmZmZmYiIiIiIiIiIiHd3d2ZmZmZmZoiIiMzMzKqqqqqqqpmZmYiIiIiIiIiIiHd3d4iIiHd3d3d3d3d3d2ZmZlVVVVVVVYiIiIiIiGZmZoiIiIiIiJmZmaqqqqqqqoiIiHd3d3d3d4iIiIiIiIiIiJmZmYiIiIiIiJmZmZmZmZmZmZmZmYiIiIiIiIiIiJmZmZmZmbu7u7u7u6qqqoiIiHd3d4iIiKqqqru7u6qqqpmZmYiIiIiIiJmZmaqqqru7u8zMzMzMzKqqqpmZmYiIiIiIiKqqqqqqqqqqqqqqqru7u5mZmYiIiIiIiJmZmbu7u6qqqru7u93d3czMzKqqqpmZmZmZmXd3d4iIiIiIiIiIiIiIiJmZmYiIiHd3d3d3d3d3d4iIiHd3d3d3d4iIiKqqqpmZmXd3d3d3d4iIiHd3d2ZmZlVVVXd3d4iIiHd3d3d3d2ZmZnd3d5mZmaqqqqqqqoiIiIiIiHd3d2ZmZnd3d3d3d3d3d1VVVXd3d3d3d3d3d3d3d3d3d3d3d4iIiJmZmaqqqpmZmXd3d4iIiHd3d2ZmZlVVVVVVVVVVVXd3d2ZmZmZmZmZmZnd3d5mZmZmZmZmZmZmZmaqqqoiIiHd3d2ZmZnd3d4iIiIiIiGZmZmZmZmZmZmZmZnd3d2ZmZnd3d4iIiJmZmaqqqqqqqqqqqoiIiHd3d4iIiHd3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZnd3d4iIiIiIiHd3d3d3d3d3d3d3d2ZmZlVVVWZmZmZmZmZmZmZmZmZmZnd3d2ZmZlVVVVVVVURERERERERERHd3d5mZmaqqqoiIiIiIiIiIiIiIiGZmZlVVVWZmZnd3d3d3d3d3d3d3d2ZmZlVVVWZmZnd3d2ZmZmZmZoiIiIiIiJmZmYiIiIiIiIiIiIiIiHd3d3d3d2ZmZnd3d4iIiHd3d3d3d3d3d3d3d3d3d2ZmZlVVVWZmZnd3d5mZmZmZmZmZmXd3d3d3d3d3d1VVVWZmZnd3d3d3d1VVVWZmZnd3d2ZmZlVVVXd3d1VVVURERERERERERFVVVURERFVVVVVVVURERERERDMzMyIiIjMzMyIiIjMzMzMzMyIiIjMzMzMzM0RERDMzM0RERFVVVVVVVVVVVTMzMzMzM1VVVXd3d3d3d4iIiGZmZmZmZlVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVURERERERERERERERERERERERFVVVWZmZlVVVVVVVWZmZlVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERERERDMzMzMzMzMzM1VVVVVVVURERFVVVURERERERDMzM0RERERERDMzMzMzM0RERFVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERCIiIjMzM1VVVVVVVURERERERERERERERDMzMzMzM0RERERERDMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzM0RERDMzMyIiIkRERGZmZkRERERERFVVVVVVVURERERERERERERERERERDMzM0RERDMzM0RERDMzMzMzM0RERERERDMzM0RERDMzMzMzM1VVVVVVVURERFVVVVVVVVVVVURERERERERERERERERERERERERERERERFVVVURERERERERERERERDMzMzMzM0RERDMzM0RERDMzMzMzMzMzMzMzM0RERFVVVVVVVURERERERFVVVVVVVVVVVURERERERERERFVVVVVVVURERDMzM1VVVVVVVVVVVTMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzM1VVVURERERERFVVVURERERERERERFVVVURERFVVVURERERERFVVVURERFVVVURERERERDMzMzMzM0RERERERERERERERERERERERFVVVVVVVURERERERERERDMzM0RERERERERERFVVVURERERERERERGZmZmZmZkRERERERERERFVVVXd3d2ZmZlVVVXd3d1VVVTMzMxERESIiIlVVVXd3d3d3d1VVVVVVVWZmZlVVVWZmZmZmZlVVVVVVVWZmZlVVVVVVVVVVVWZmZlVVVURERDMzM0RERERERERERFVVVVVVVWZmZoiIiJmZmYiIiHd3d3d3d2ZmZlVVVTMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERFVVVURERFVVVURERERERERERERERDMzMzMzM0RERDMzM0RERERERDMzMzMzMzMzMzMzMyIiIiIiIiIiIjMzMyIiIiIiIjMzMyIiIjMzMzMzMzMzM0RERFVVVVVVVVVVVURERERERERERERERERERERERFVVVVVVVVVVVURERERERERERERERERERERERERERGZmZmZmZkRERFVVVURERERERERERFVVVWZmZmZmZlVVVURERERERFVVVVVVVXd3d2ZmZnd3d3d3d4iIiIiIiJmZmaqqqqqqqmZmZkRERCIiIlVVVaqqqpmZmXd3d1VVVURERDMzMzMzM0RERERERERERFVVVURERERERFVVVXd3d3d3d1VVVURERERERFVVVWZmZlVVVURERERERFVVVXd3d2ZmZmZmZnd3d4iIiIiIiFVVVVVVVVVVVVVVVURERFVVVVVVVVVVVXd3d3d3d3d3d2ZmZnd3d4iIiFVVVVVVVVVVVVVVVXd3d5mZmXd3d3d3d7u7u6qqqmZmZmZmZnd3d2ZmZmZmZmZmZlVVVVVVVVVVVXd3d4iIiGZmZlVVVVVVVWZmZkRERERERGZmZnd3d2ZmZlVVVURERFVVVVVVVVVVVYiIiJmZmYiIiFVVVURERGZmZlVVVURERERERERERERERFVVVVVVVWZmZmZmZmZmZkRERFVVVVVVVURERFVVVURERERERFVVVVVVVVVVVWZmZnd3d1VVVVVVVWZmZoiIiHd3d2ZmZmZmZmZmZoiIiIiIiGZmZlVVVVVVVVVVVVVVVXd3d3d3d3d3d1VVVVVVVURERGZmZmZmZnd3d6qqqt3d3bu7u4iIiFVVVVVVVYiIiHd3d3d3d2ZmZkRERDMzM0RERERERERERERERFVVVURERERERFVVVWZmZmZmZmZmZmZmZoiIiLu7u+7u7v///////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3d3d3MzMzMzMy7u7u7u7vMzMzMzMzMzMzMzMzMzMzMzMzd3d3d3d3MzMzd3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7d3d3u7u7d3d3MzMy7u7u7u7u7u7uqqqqZmZmqqqqZmZmZmZmZmZmIiIiIiIiZmZmZmZmIiIiIiIiIiIh3d3d3d3eIiIiIiIiIiIh3d3eIiIiIiIh3d3eIiIiIiIiIiIh3d3d3d3eIiIiIiIh3d3d3d3eIiIh3d3eIiIiIiIiIiIh3d3eIiIiIiIh3d3d3d3eIiIiIiIiIiIiZmZmZmZmIiIiIiIiIiIh3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIiIiIiIiIh3d3d3d3d3d3d3d3eIiIh3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVEREREREREREREREREREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNERERVVVVERERERERERERERERERERVVVV3d3dmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZ3d3dVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVV3d3eZmZm7u7uZmZl3d3eIiIiqqqqqqqqIiIiIiIiIiIhmZmZVVVVVVVVERERVVVVVVVVERERVVVVmZmZVVVVEREREREQzMzNVVVWIiIjMzMzd3d3MzMzd3d3MzMzMzMy7u7u7u7uqqqqZmZmqqqqZmZmIiIiIiIiIiIiIiIiIiIh3d3eIiIi7u7vMzMyZmZmZmZl3d3dmZmZ3d3eIiIiZmZl3d3d3d3d3d3dmZmZmZmZmZmaIiIh3d3d3d3eIiIiIiIiIiIiqqqqqqqqZmZl3d3eIiIiIiIiZmZmZmZmZmZmIiIiIiIiZmZmZmZmqqqqqqqqZmZmIiIiIiIiZmZmZmZmZmZmZmZmZmZl3d3eIiIiZmZmqqqq7u7uqqqqZmZmIiIiZmZm7u7vMzMy7u7u7u7uqqqqZmZmqqqqIiIh3d3eZmZmqqqqqqqqqqqqZmZmIiIiIiIiZmZmqqqq7u7u7u7vMzMzMzMy7u7uIiIh3d3eIiIh3d3d3d3eIiIiZmZmZmZmIiIh3d3d3d3d3d3eIiIiIiIiIiIiZmZmqqqqqqqqIiIiIiIiIiIh3d3dVVVVmZmZ3d3d3d3dmZmZmZmaIiIh3d3eIiIiqqqqqqqqZmZmIiIiIiIh3d3dmZmZmZmaIiIiIiIhVVVVmZmZ3d3d3d3d3d3d3d3dmZmaIiIiqqqqqqqqIiIhmZmZ3d3d3d3dVVVV3d3dmZmZmZmZ3d3dmZmZVVVVmZmZ3d3eZmZmZmZmZmZmZmZmZmZmZmZmIiIh3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3dmZmZ3d3d3d3eIiIiZmZmqqqqqqqqqqqqIiIiIiIh3d3d3d3d3d3d3d3dmZmZ3d3d3d3dmZmZ3d3dmZmaIiIiIiIh3d3d3d3d3d3dmZmZmZmZmZmZmZmZVVVVmZmZmZmZVVVV3d3dmZmZmZmZmZmZVVVUzMzNVVVWIiIiqqqqZmZmIiIiZmZmZmZl3d3dmZmZmZmZmZmZ3d3d3d3d3d3d3d3dmZmZVVVVmZmZVVVVVVVVmZmaIiIiZmZmZmZmZmZmIiIiZmZmIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dERERVVVV3d3eZmZmIiIiIiIh3d3dmZmZmZmZ3d3d3d3d3d3dmZmZVVVVVVVVmZmZmZmZVVVV3d3dmZmZERERERERERERVVVVERERERERVVVVEREQzMzMiIiIiIiIzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzNERER3d3d3d3d3d3eIiIh3d3dVVVVmZmZVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVEREREREREREQzMzNERERVVVVmZmZVVVVmZmZVVVVVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVEREREREREREQzMzMzMzMzMzNVVVVERERVVVVmZmZVVVVEREQzMzMzMzMzMzNEREQzMzNERERVVVUzMzMzMzMzMzMzMzNEREQzMzMiIiJEREREREQzMzNERERVVVVVVVVVVVVEREREREQzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzNEREQzMzMzMzNERERmZmZERERERERERERVVVVVVVVEREREREREREREREREREREREQzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzNERERERERVVVVERERERERVVVVVVVVVVVVVVVVERERERERERERERERERERERERVVVVEREREREREREQzMzNEREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzNEREQzMzNVVVVERERERERERERVVVVERERVVVVERERERERERERVVVVEREQzMzNERERVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzNERERERERERERERERERERVVVVERERERERERERVVVVERERERERERERERERVVVVEREREREREREREREREREREREQzMzNERERERERERERERERVVVVERERVVVVEREREREREREREREQzMzNERERERERVVVVVVVVVVVVVVVUzMzMzMzNVVVV3d3eIiIhVVVVEREREREREREQiIiIiIiIiIiJERER3d3d3d3dmZmZVVVVmZmZmZmZmZmZVVVVVVVVVVVVmZmZERERVVVVVVVVVVVVVVVVEREQzMzNERERERERVVVV3d3dmZmZVVVWZmZmqqqqIiIh3d3d3d3d3d3dVVVVEREREREQzMzMzMzMiIiIiIiIzMzMzMzNERERERERERERERERVVVVVVVVVVVVEREREREREREREREQzMzMzMzNERERVVVVEREREREREREREREQzMzMzMzMzMzMiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIiIiJERERVVVVmZmZVVVUzMzNERERERERVVVVERERVVVVERERVVVVVVVVERERVVVVEREQzMzNVVVVVVVUzMzNERERVVVVVVVVERERERERERERERERERERVVVV3d3dVVVVVVVVERERERERVVVVVVVVmZmZmZmZ3d3d3d3d3d3eIiIiZmZmqqqqZmZlVVVVEREQiIiJERES7u7uZmZl3d3dERERERERERERERERERERERERVVVVVVVVERERERERVVVVVVVVmZmZVVVVERERERERVVVVVVVVmZmZVVVVVVVVmZmZmZmZVVVVVVVVmZmaIiIiIiIhmZmZERERVVVVVVVVVVVVVVVVVVVVVVVV3d3d3d3dVVVVVVVVVVVVVVVVVVVVVVVVVVVV3d3d3d3eZmZmZmZmZmZnMzMyZmZlVVVVmZmZmZmZmZmZERERERERERERVVVVmZmZmZmZmZmZVVVVVVVVVVVVmZmZERERERERmZmZmZmZERERERERERERVVVVERERERER3d3e7u7uIiIhVVVVVVVVmZmZVVVVERERERERERERERERERERVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVERERVVVVVVVV3d3dmZmZVVVV3d3eIiIh3d3dmZmZ3d3d3d3eIiIiZmZlmZmZERERERERVVVVmZmaIiIiIiIh3d3dVVVVVVVVVVVVmZmZ3d3eZmZmqqqrMzMyZmZlmZmZmZmZmZmaIiIh3d3dVVVVERERERERERERERERERERVVVVVVVVERERERERVVVVmZmaIiIhmZmZmZmaZmZm7u7vd3d3///////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7uzMzMu7u7u7u7u7u7zMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d7u7u7u7u3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMu7u7u7u7qqqqmZmZmZmZmZmZqqqqmZmZmZmZiIiId3d3iIiIiIiId3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmd3d3d3d3d3d3ZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3iIiIZmZmVVVVZmZmZmZmZmZmd3d3d3d3ZmZmZmZmVVVVZmZmZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3iIiIiIiImZmZmZmZiIiIiIiIiIiId3d3d3d3iIiId3d3iIiId3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmd3d3d3d3ZmZmVVVVVVVVZmZmZmZmZmZmVVVVZmZmiIiImZmZu7u7qqqqiIiIiIiIqqqqu7u7iIiId3d3d3d3d3d3VVVVREREREREREREVVVVREREVVVVREREVVVVREREMzMzREREZmZmmZmZzMzM3d3d3d3dzMzMzMzMqqqqu7u7qqqqqqqqu7u7u7u7qqqqd3d3d3d3iIiIqqqqmZmZmZmZiIiIqqqqu7u7qqqqiIiId3d3d3d3d3d3mZmZiIiIiIiId3d3d3d3iIiIiIiIiIiImZmZiIiId3d3d3d3ZmZmZmZmmZmZu7u7mZmZiIiIiIiImZmZiIiId3d3iIiIiIiId3d3iIiImZmZu7u7mZmZiIiIiIiImZmZmZmZd3d3ZmZmqqqqqqqqmZmZmZmZqqqqqqqqqqqqmZmZiIiImZmZzMzM3d3d3d3dzMzMu7u7u7u7u7u7mZmZiIiIZmZmiIiIqqqqmZmZmZmZmZmZiIiImZmZqqqqqqqqu7u7u7u7u7u7qqqqqqqqiIiIiIiId3d3iIiId3d3iIiIiIiIiIiIiIiId3d3iIiImZmZiIiImZmZmZmZqqqqmZmZmZmZmZmZiIiIiIiId3d3VVVVZmZmd3d3ZmZmZmZmd3d3d3d3iIiIqqqqu7u7qqqqmZmZd3d3mZmZd3d3d3d3ZmZmiIiImZmZd3d3d3d3iIiId3d3ZmZmZmZmiIiImZmZmZmZqqqqiIiIiIiImZmZd3d3ZmZmd3d3d3d3d3d3ZmZmZmZmZmZmd3d3iIiIiIiIiIiImZmZqqqqmZmZiIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmd3d3d3d3d3d3iIiImZmZmZmZqqqqqqqqmZmZd3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmd3d3ZmZmd3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3VVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmZmZmREREVVVViIiImZmZmZmZmZmZmZmZmZmZiIiIiIiId3d3ZmZmd3d3d3d3d3d3d3d3d3d3ZmZmZmZmREREREREVVVViIiImZmZqqqqqqqqiIiIiIiIiIiIiIiImZmZiIiId3d3d3d3d3d3iIiIiIiId3d3d3d3VVVVREREVVVVd3d3iIiImZmZiIiId3d3ZmZmd3d3d3d3d3d3mZmZd3d3ZmZmZmZmd3d3ZmZmZmZmZmZmZmZmREREREREREREVVVVREREREREVVVVMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzREREREREMzMzREREVVVVd3d3iIiIZmZmd3d3ZmZmZmZmZmZmVVVVREREVVVVREREVVVVVVVVVVVVVVVVREREREREREREREREREREZmZmZmZmVVVVVVVVZmZmREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREREREMzMzREREREREREREVVVVZmZmVVVVREREREREREREMzMzREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREMzMzREREVVVVREREREREVVVVREREMzMzMzMzREREMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzREREMzMzMzMzREREVVVVREREREREREREVVVVREREREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREVVVVREREVVVVVVVVREREREREVVVVREREREREREREVVVVREREMzMzREREREREREREREREREREMzMzREREMzMzMzMzMzMzREREMzMzREREREREREREVVVVREREREREREREREREREREVVVVVVVVREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiREREREREREREREREREREREREREREVVVVREREREREVVVVREREREREREREREREREREREREMzMzREREREREMzMzMzMzMzMzREREREREREREVVVVREREREREREREREREREREREREREREREREREREREREVVVVZmZmREREREREREREd3d3iIiIZmZmREREREREMzMzMzMzIiIiERERIiIiMzMzd3d3d3d3d3d3ZmZmVVVVZmZmd3d3VVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVREREMzMzREREMzMzREREVVVVVVVVZmZmiIiImZmZmZmZd3d3iIiId3d3ZmZmREREMzMzMzMzREREMzMzMzMzMzMzMzMzREREMzMzREREVVVVREREVVVVREREREREMzMzMzMzMzMzMzMzMzMzVVVVZmZmVVVVVVVVVVVVREREMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzIiIiIiIiREREVVVVREREREREMzMzMzMzMzMzMzMzVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREREREREREREREREREREREREREREREREREREREMzMzREREZmZmd3d3VVVVREREREREREREVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3qqqqu7u7mZmZZmZmMzMzIiIiVVVVqqqqmZmZZmZmVVVVREREREREMzMzREREREREVVVVREREREREREREVVVVVVVVVVVVVVVVREREVVVVVVVVREREVVVVZmZmZmZmVVVVVVVVREREREREVVVVZmZmd3d3ZmZmREREREREZmZmVVVVVVVVREREVVVVZmZmd3d3VVVVREREVVVVVVVVZmZmVVVVd3d3mZmZiIiIqqqqzMzMmZmZu7u7iIiIZmZmZmZmVVVVREREVVVVVVVVVVVVd3d3ZmZmVVVVREREZmZmVVVVREREVVVVREREREREREREREREREREREREREREVVVVVVVVREREZmZmu7u7mZmZVVVVZmZmVVVVREREMzMzMzMzMzMzREREREREZmZmd3d3VVVVVVVVd3d3ZmZmVVVVVVVVVVVVREREVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmd3d3mZmZiIiIZmZmd3d3d3d3iIiId3d3ZmZmREREREREVVVVZmZmiIiIiIiId3d3VVVVVVVVVVVVd3d3mZmZqqqqu7u7mZmZd3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREREREVVVVZmZmREREVVVVVVVVZmZmd3d3d3d3ZmZmiIiIzMzM////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////+7u7szMzLu7u7u7u8zMzN3d3d3d3d3d3e7u7t3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3czMzMzMzN3d3czMzN3d3czMzN3d3d3d3d3d3d3d3e7u7t3d3d3d3e7u7t3d3d3d3d3d3czMzMzMzLu7u7u7u6qqqpmZmZmZmZmZmXd3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVURERERERERERFVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZnd3d2ZmZmZmZnd3d4iIiGZmZlVVVURERFVVVVVVVWZmZmZmZmZmZlVVVWZmZlVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d4iIiIiIiIiIiJmZmZmZmYiIiIiIiJmZmZmZmYiIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d2ZmZmZmZnd3d3d3d2ZmZlVVVWZmZmZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVXd3d3d3d2ZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVYiIiJmZmaqqqnd3d3d3d4iIiJmZmaqqqpmZmWZmZnd3d3d3d2ZmZkRERERERFVVVURERFVVVVVVVVVVVVVVVVVVVURERFVVVYiIiLu7u8zMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u6qqqqqqqqqqqoiIiHd3d4iIiJmZmaqqqqqqqoiIiGZmZoiIiKqqqpmZmZmZmYiIiHd3d3d3d3d3d3d3d2ZmZoiIiIiIiIiIiKqqqru7u7u7u4iIiGZmZmZmZlVVVXd3d5mZmaqqqqqqqoiIiIiIiIiIiHd3d3d3d3d3d3d3d4iIiJmZmaqqqqqqqpmZmWZmZmZmZpmZmYiIiFVVVVVVVYiIiKqqqpmZmaqqqpmZmaqqqpmZmXd3d5mZmd3d3d3d3d3d3bu7u7u7u7u7u6qqqpmZmYiIiHd3d3d3d4iIiJmZmYiIiIiIiIiIiJmZmaqqqqqqqqqqqru7u6qqqqqqqpmZmaqqqpmZmYiIiHd3d6qqqpmZmXd3d3d3d3d3d3d3d3d3d5mZmYiIiIiIiKqqqru7u5mZmYiIiIiIiHd3d3d3d4iIiHd3d3d3d3d3d3d3d2ZmZmZmZnd3d3d3d6qqqru7u6qqqoiIiIiIiIiIiJmZmYiIiHd3d2ZmZoiIiJmZmXd3d2ZmZmZmZmZmZmZmZnd3d5mZmbu7u6qqqqqqqpmZmZmZmYiIiHd3d2ZmZnd3d4iIiHd3d2ZmZmZmZnd3d4iIiIiIiIiIiJmZmZmZmaqqqoiIiIiIiIiIiIiIiIiIiGZmZmZmZnd3d3d3d1VVVWZmZnd3d2ZmZnd3d4iIiJmZmZmZmbu7u6qqqpmZmYiIiHd3d3d3d2ZmZmZmZlVVVWZmZmZmZmZmZmZmZnd3d4iIiHd3d3d3d3d3d3d3d3d3d4iIiHd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmXd3d3d3d4iIiHd3d3d3d2ZmZnd3d2ZmZmZmZnd3d4iIiHd3d3d3d2ZmZkRERERERGZmZoiIiIiIiJmZmZmZmYiIiIiIiIiIiJmZmaqqqpmZmYiIiHd3d4iIiJmZmYiIiHd3d2ZmZkRERERERGZmZoiIiIiIiIiIiJmZmZmZmXd3d2ZmZmZmZoiIiIiIiIiIiGZmZlVVVWZmZlVVVWZmZmZmZlVVVVVVVURERERERDMzMzMzM0RERERERERERDMzMzMzMyIiIiIiIjMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzM0RERERERERERERERGZmZmZmZmZmZnd3d2ZmZlVVVVVVVVVVVURERERERERERERERERERERERERERERERERERERERERERFVVVWZmZmZmZkRERFVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVTMzMzMzM1VVVURERERERERERERERERERERERERERFVVVURERERERERERERERERERERERERERERERDMzMzMzM0RERERERDMzMzMzM0RERERERERERERERERERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMyIiIjMzM0RERFVVVTMzM0RERERERERERFVVVURERDMzMzMzMzMzM0RERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERERERFVVVVVVVURERERERERERERERERERDMzMzMzM0RERERERERERDMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzM0RERDMzMzMzM0RERERERERERFVVVURERERERFVVVVVVVURERERERERERDMzMzMzM0RERERERERERDMzM0RERERERERERERERDMzMzMzMzMzMyIiIjMzMzMzM0RERERERERERERERERERERERFVVVURERERERERERFVVVURERERERERERDMzMzMzM0RERERERDMzMzMzM0RERERERERERFVVVVVVVURERERERERERDMzMzMzMzMzM0RERERERFVVVVVVVURERFVVVVVVVVVVVVVVVWZmZnd3d2ZmZkRERERERDMzMzMzMzMzMyIiIiIiIhERETMzM1VVVYiIiIiIiGZmZmZmZmZmZmZmZlVVVURERERERERERFVVVVVVVWZmZlVVVURERDMzMzMzM0RERDMzM0RERERERERERGZmZnd3d5mZmZmZmXd3d2ZmZnd3d2ZmZlVVVTMzMzMzM0RERDMzMzMzM0RERERERERERDMzM0RERERERERERERERERERERERDMzMzMzMzMzMyIiIkRERHd3d2ZmZlVVVVVVVURERERERERERDMzMzMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzM0RERDMzMzMzM0RERFVVVVVVVVVVVURERERERFVVVURERDMzM0RERFVVVURERERERERERDMzMzMzM0RERDMzM0RERERERFVVVVVVVWZmZlVVVURERERERGZmZnd3d2ZmZlVVVXd3d2ZmZmZmZnd3d6qqqt3d3aqqqmZmZkRERCIiIkRERJmZmXd3d1VVVVVVVURERERERERERERERERERERERERERERERERERFVVVXd3d4iIiHd3d1VVVVVVVWZmZkRERERERFVVVVVVVVVVVURERERERERERERERFVVVVVVVVVVVURERFVVVVVVVVVVVVVVVURERERERHd3d3d3d2ZmZmZmZmZmZmZmZnd3d3d3d5mZmbu7u6qqqru7u8zMzJmZmZmZmYiIiFVVVURERFVVVVVVVWZmZmZmZmZmZlVVVURERERERFVVVXd3d2ZmZkRERERERFVVVURERERERERERERERERERERERFVVVVVVVURERHd3d7u7u4iIiFVVVVVVVTMzMzMzMyIiIjMzMzMzMzMzM0RERGZmZnd3d0RERFVVVWZmZmZmZmZmZlVVVURERFVVVURERFVVVURERFVVVVVVVVVVVXd3d4iIiJmZmaqqqoiIiHd3d2ZmZnd3d3d3d2ZmZlVVVURERFVVVWZmZnd3d3d3d4iIiGZmZmZmZmZmZnd3d4iIiLu7u93d3bu7u4iIiGZmZnd3d3d3d1VVVVVVVVVVVWZmZlVVVVVVVURERERERFVVVVVVVWZmZmZmZnd3d2ZmZmZmZlVVVXd3d7u7u+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////u7u7////u7u7MzMzMzMzd3d3u7u7d3d3d3d3MzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3d3d3u7u7d3d3u7u7d3d3u7u7d3d3d3d3u7u7d3d3d3d3d3d3d3d3MzMzd3d3d3d3MzMzMzMzMzMzMzMy7u7vMzMy7u7u7u7uqqqqZmZmZmZmIiIiIiIh3d3dmZmZmZmZmZmZVVVVmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZ3d3d3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3eIiIiIiIiIiIiIiIiZmZmIiIiIiIiIiIh3d3dmZmZ3d3d3d3eIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3eIiIh3d3d3d3eIiIh3d3d3d3eIiIh3d3eIiIiIiIiIiIiZmZmZmZmIiIiIiIiZmZmIiIiIiIiIiIiIiIh3d3eIiIiIiIiIiIh3d3d3d3d3d3dmZmZmZmZmZmZVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERERERVVVVERERVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZVVVVmZmaIiIiqqqqqqqqIiIh3d3eIiIiqqqqZmZl3d3dmZmZ3d3eZmZl3d3dVVVVERERERERVVVVmZmZmZmZVVVVVVVVVVVVVVVVmZmaZmZm7u7u7u7u7u7vd3d3MzMzd3d27u7u7u7u7u7uqqqqZmZmqqqp3d3eZmZm7u7u7u7uqqqqZmZl3d3dmZmZmZmaIiIiqqqqZmZl3d3d3d3dVVVVmZmZmZmZmZmZmZmZ3d3eqqqqqqqqZmZmIiIh3d3dmZmZVVVVVVVVmZmZ3d3eZmZmZmZmIiIh3d3d3d3dmZmZ3d3eIiIiIiIiZmZmqqqqqqqqqqqqZmZmIiIhmZmZ3d3d3d3dVVVVVVVV3d3eIiIiZmZmqqqqqqqqZmZmIiIh3d3eqqqrd3d3d3d3MzMzMzMy7u7u7u7uZmZmIiIh3d3eIiIiIiIiZmZmIiIiIiIh3d3eIiIiIiIiqqqqqqqqqqqq7u7uqqqqZmZmqqqqqqqqqqqqIiIiIiIiqqqqZmZmIiIhmZmZmZmZ3d3eIiIh3d3d3d3eIiIiqqqqqqqqIiIh3d3eIiIh3d3d3d3d3d3d3d3eIiIh3d3dmZmZmZmZmZmZmZmaIiIiqqqq7u7uqqqqZmZmIiIiZmZmZmZmIiIh3d3dVVVV3d3eZmZmIiIhmZmZERERVVVVmZmaIiIiqqqqZmZmqqqqqqqqZmZmIiIiIiIh3d3d3d3d3d3dmZmZ3d3dmZmZmZmZVVVVmZmaIiIiIiIiZmZmZmZmZmZmZmZmIiIiIiIiIiIh3d3d3d3dmZmZ3d3d3d3dmZmZERERVVVV3d3eIiIiZmZmZmZmZmZmZmZmIiIh3d3eZmZmIiIiIiIhmZmZmZmZVVVVmZmZmZmZVVVVmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3eIiIhmZmZmZmZmZmZmZmZmZmZmZmZ3d3dVVVVVVVVVVVVVVVV3d3d3d3eZmZmIiIh3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3eIiIiZmZl3d3d3d3dmZmZVVVVERERVVVV3d3eIiIiZmZmZmZmqqqqZmZmZmZmIiIiIiIiZmZmZmZl3d3eIiIiIiIh3d3dmZmZVVVVVVVVERERmZmaIiIiIiIiIiIiZmZmIiIh3d3dmZmZ3d3dmZmZ3d3d3d3dmZmZVVVVmZmZmZmZVVVVmZmZVVVVVVVUzMzMzMzNEREREREQzMzNERERVVVVEREQzMzMiIiIzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMzMzNVVVVEREQzMzNERERERERmZmZ3d3d3d3dmZmZmZmZVVVVVVVVVVVVEREQzMzNERERERERERERERERERERERERERERERERVVVVVVVVVVVVVVVVERERVVVVVVVVERERVVVVERERVVVVERERERERERERVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVERERERERERERERERERERERERERERERERERERERERVVVVVVVVERERERERVVVVVVVVEREREREREREREREREREREREREREREREQzMzNERERERERVVVVEREREREREREREREQzMzNEREREREQzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzNEREQzMzMiIiJERERVVVVERERERERERERERERERERERERERERVVVVEREREREREREREREQzMzNEREREREQzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzNEREREREREREREREREREREREREREQzMzNEREQzMzMzMzNEREREREQzMzNEREREREREREREREREREREREQzMzMzMzMiIiIzMzMzMzMzMzNERERERERERERVVVVVVVVERERERERERERERERERERERERVVVVEREREREREREREREREREREREREREREREREREREREREREQzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREREREREREREREREREREREREREREREQzMzNEREQzMzNEREREREQzMzMzMzNERERERERERERVVVVVVVVERERERERERERERERERERERERERERERERERERERERVVVVVVVVVVVVmZmZVVVVmZmZVVVVmZmZEREQzMzMzMzMiIiIzMzMzMzMiIiIREREiIiJVVVV3d3d3d3dmZmZmZmZmZmZmZmZEREREREQzMzNERERVVVVVVVVVVVVVVVVEREREREQzMzNEREQzMzMzMzNERERERERVVVVmZmaZmZmqqqqIiIhmZmZmZmZ3d3dVVVVERERERERERERERERERERVVVVVVVVEREQzMzNEREREREREREREREREREREREREREREREQzMzMzMzN3d3eIiIhmZmZEREREREREREREREREREREREQzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzNERERVVVVVVVVVVVVEREREREREREQzMzNERERVVVVEREREREREREREREREREREREREREQzMzNERERERERVVVVVVVVVVVVVVVVERERVVVV3d3dmZmZmZmZmZmZmZmZVVVVVVVWIiIjMzMzMzMx3d3dEREQiIiIzMzN3d3eIiIhmZmZERERERERVVVVERERERERERERERERERERERERVVVV3d3eZmZm7u7uqqqpmZmZVVVVERERVVVVERERERERVVVVmZmZVVVVERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVERER3d3dmZmZmZmZmZmZmZmZmZmZ3d3d3d3eZmZmqqqqqqqq7u7uqqqp3d3eZmZl3d3dVVVVVVVVVVVVVVVVmZmZVVVVERERVVVVERERERERVVVV3d3dmZmZEREREREREREQzMzMzMzNERERERERERERVVVVVVVVmZmZmZmZmZmaIiIh3d3dVVVVERERERERERERERERVVVVEREQzMzMzMzNVVVVmZmZmZmZVVVVERERERERmZmZVVVVVVVVERERVVVVERERERERVVVVVVVVVVVV3d3d3d3eqqqqZmZl3d3dmZmZmZmaIiIh3d3dVVVVERERERERVVVVVVVVmZmaIiIh3d3dmZmZmZmZmZmaZmZm7u7vMzMy7u7uZmZl3d3eIiIh3d3dERERERERVVVVVVVVmZmZVVVVVVVVERERVVVVmZmZ3d3eIiIh3d3dmZmZVVVVVVVVmZmaIiIiqqqrd3d3u7u7////u7u7u7u7u7u7////u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7////u7u7///////////////////////////////////////////////////////8A////////////////////7u7u////////////////////////////////////////7u7u////////////7u7u////////7u7u////////////////////////7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3dzMzMzMzM3d3d3d3d3d3d7u7u3d3d7u7u3d3d3d3d7u7u3d3d7u7u3d3d3d3dzMzMzMzMzMzMu7u7u7u7u7u7u7u7u7u7u7u7qqqqu7u7u7u7u7u7u7u7u7u7u7u7zMzMu7u7zMzMu7u7u7u7qqqqmZmZmZmZqqqqmZmZmZmZmZmZmZmZiIiImZmZmZmZiIiIiIiImZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZiIiIiIiImZmZmZmZmZmZmZmZmZmZmZmZqqqqmZmZmZmZqqqqmZmZmZmZiIiImZmZqqqqqqqqqqqqmZmZmZmZmZmZmZmZiIiIiIiIiIiImZmZiIiImZmZiIiId3d3iIiId3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmd3d3d3d3ZmZmd3d3d3d3ZmZmd3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREREREREREREREREREMzMzMzMzREREREREREREMzMzMzMzMzMzREREREREREREREREREREREREVVVVVVVVVVVVREREVVVVZmZmZmZmiIiIqqqqqqqqmZmZiIiIiIiIiIiIiIiId3d3ZmZmd3d3mZmZZmZmVVVVREREVVVVREREVVVVZmZmZmZmZmZmVVVVVVVVVVVVZmZmiIiIqqqqu7u7zMzMzMzMzMzMqqqqqqqqzMzMqqqqmZmZmZmZmZmZmZmZu7u7qqqqiIiIZmZmZmZmd3d3d3d3d3d3mZmZmZmZiIiIZmZmVVVVZmZmZmZmd3d3ZmZmmZmZu7u7mZmZZmZmZmZmZmZmZmZmVVVVZmZmZmZmd3d3iIiIiIiId3d3iIiId3d3d3d3iIiIiIiImZmZu7u7qqqqqqqqmZmZiIiIiIiId3d3ZmZmZmZmZmZmVVVVZmZmmZmZqqqqmZmZmZmZiIiId3d3mZmZzMzM7u7uzMzMzMzMu7u7qqqqqqqqqqqqiIiIZmZmiIiImZmZiIiIiIiId3d3d3d3d3d3iIiIqqqqqqqqqqqqu7u7qqqqqqqqqqqqmZmZmZmZiIiIiIiImZmZmZmZiIiIZmZmd3d3d3d3d3d3d3d3d3d3mZmZqqqqmZmZiIiId3d3d3d3iIiIiIiId3d3iIiIiIiId3d3ZmZmZmZmZmZmZmZmqqqqu7u7u7u7qqqqqqqqmZmZqqqqmZmZiIiIZmZmVVVVZmZmiIiIiIiIZmZmVVVVd3d3iIiImZmZqqqqmZmZmZmZmZmZiIiIiIiIiIiId3d3d3d3ZmZmZmZmZmZmd3d3ZmZmVVVVZmZmiIiImZmZqqqqmZmZmZmZmZmZd3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3ZmZmREREVVVVd3d3mZmZmZmZmZmZmZmZmZmZiIiIiIiImZmZiIiIiIiIiIiId3d3ZmZmZmZmVVVVZmZmVVVVd3d3d3d3d3d3d3d3iIiId3d3d3d3iIiId3d3d3d3ZmZmd3d3d3d3d3d3d3d3ZmZmVVVVZmZmVVVVZmZmd3d3iIiIiIiIiIiId3d3iIiIiIiIiIiIiIiId3d3d3d3iIiId3d3d3d3iIiId3d3VVVVVVVVREREREREZmZmd3d3mZmZiIiIqqqqqqqqiIiIiIiIiIiIiIiImZmZmZmZiIiId3d3d3d3ZmZmZmZmVVVVVVVVVVVVd3d3mZmZmZmZmZmZmZmZmZmZd3d3ZmZmZmZmZmZmVVVVZmZmZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREREREREREMzMzMzMzVVVVREREREREMzMzIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzIiIiMzMzMzMzREREREREREREVVVVd3d3d3d3ZmZmd3d3ZmZmVVVVVVVVVVVVVVVVREREVVVVREREMzMzMzMzREREREREREREVVVVREREREREVVVVREREVVVVVVVVREREVVVVVVVVREREVVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREMzMzMzMzREREMzMzREREREREVVVVZmZmVVVVVVVVZmZmVVVVVVVVVVVVREREVVVVREREREREREREREREREREMzMzREREVVVVREREZmZmVVVVREREREREREREMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzREREIiIiMzMzMzMzVVVVREREMzMzREREREREMzMzREREREREVVVVVVVVREREMzMzMzMzREREREREMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVVVVVREREVVVVREREREREREREREREREREMzMzMzMzMzMzREREMzMzREREREREREREMzMzREREMzMzREREMzMzMzMzMzMzIiIiMzMzMzMzREREREREREREREREREREREREREREMzMzMzMzREREREREREREREREREREREREREREREREREREREREREREREREREREMzMzIiIiMzMzMzMzMzMzREREREREREREREREREREREREREREREREMzMzREREMzMzREREMzMzMzMzREREREREREREMzMzREREMzMzREREREREVVVVVVVVVVVVREREREREREREMzMzREREREREREREREREREREVVVVVVVVZmZmiIiIZmZmZmZmVVVVREREVVVVREREMzMzMzMzMzMzMzMzIiIiMzMzREREVVVVZmZmVVVVZmZmZmZmZmZmVVVVREREMzMzREREREREREREVVVVREREREREREREREREREREREREMzMzREREMzMzMzMzREREZmZmd3d3mZmZmZmZd3d3d3d3ZmZmVVVVVVVVVVVVREREREREVVVVVVVVVVVVREREREREMzMzREREREREREREVVVVREREREREMzMzMzMzVVVVqqqqiIiIVVVVMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiREREREREMzMzIiIiMzMzMzMzREREREREREREREREREREMzMzVVVVVVVVREREVVVVREREREREMzMzREREVVVVREREMzMzREREREREMzMzREREREREREREREREVVVVREREREREVVVVREREVVVVVVVVd3d3ZmZmVVVVZmZmZmZmZmZmZmZmmZmZ3d3dzMzMd3d3REREIiIiMzMzd3d3iIiIZmZmVVVVREREVVVVREREREREREREVVVVREREREREZmZmiIiImZmZmZmZmZmZd3d3VVVVREREVVVVREREREREVVVVVVVVVVVVVVVVREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVREREREREZmZmZmZmVVVVVVVVVVVVVVVVZmZmiIiImZmZiIiImZmZu7u7iIiId3d3d3d3ZmZmREREVVVVREREREREVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmVVVVREREMzMzMzMzREREMzMzREREREREVVVVVVVVZmZmZmZmZmZmZmZmd3d3d3d3VVVVREREVVVVREREVVVVVVVVVVVVREREREREREREVVVVZmZmVVVVREREREREZmZmd3d3ZmZmVVVVREREVVVVVVVVREREREREVVVVZmZmd3d3qqqqqqqqZmZmVVVVZmZmd3d3d3d3REREREREVVVVVVVVVVVVd3d3mZmZd3d3d3d3d3d3mZmZzMzMzMzMmZmZiIiId3d3iIiId3d3REREREREVVVVZmZmVVVVVVVVVVVVVVVVREREVVVVd3d3d3d3d3d3ZmZmREREREREZmZmiIiIiIiIiIiIqqqqu7u7u7u7mZmZiIiIqqqqu7u7u7u7u7u7u7u7u7u7qqqqu7u7zMzMu7u7u7u7zMzMzMzM7u7u7u7u////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7u7u7u7u7u7u7u7u7t3d3d3d3e7u7t3d3d3d3d3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3d3d3czMzMzMzMzMzLu7u8zMzMzMzMzMzLu7u6qqqpmZmYiIiJmZmZmZmaqqqqqqqqqqqru7u7u7u8zMzMzMzMzMzMzMzN3d3czMzN3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u7u7u6qqqqqqqqqqqpmZmZmZmaqqqqqqqqqqqru7u6qqqpmZmZmZmaqqqqqqqqqqqqqqqqqqqpmZmaqqqpmZmYiIiIiIiIiIiIiIiIiIiIiIiJmZmYiIiIiIiJmZmYiIiHd3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERERERERERERERERERERERERERERERERERERERERERERERERERERERFVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERDMzM0RERDMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzM0RERERERERERDMzM0RERERERFVVVURERERERGZmZmZmZmZmZlVVVVVVVURERERERFVVVWZmZnd3d3d3d3d3d5mZmZmZmXd3d3d3d4iIiHd3d2ZmZmZmZnd3d5mZmXd3d1VVVVVVVWZmZmZmZmZmZnd3d3d3d3d3d1VVVURERFVVVURERGZmZnd3d5mZmaqqqqqqqru7u7u7u7u7u7u7u6qqqpmZmaqqqru7u6qqqqqqqoiIiHd3d2ZmZmZmZmZmZoiIiIiIiHd3d3d3d4iIiHd3d3d3d2ZmZlVVVWZmZoiIiKqqqpmZmYiIiGZmZnd3d2ZmZlVVVWZmZmZmZlVVVXd3d4iIiIiIiHd3d4iIiIiIiHd3d5mZmYiIiKqqqru7u7u7u4iIiIiIiIiIiIiIiHd3d2ZmZnd3d2ZmZmZmZnd3d6qqqqqqqpmZmZmZmYiIiHd3d7u7u93d3czMzKqqqqqqqpmZmZmZmaqqqqqqqoiIiGZmZnd3d5mZmZmZmZmZmXd3d3d3d2ZmZpmZmbu7u6qqqpmZmaqqqru7u7u7u7u7u5mZmZmZmYiIiIiIiIiIiJmZmZmZmXd3d2ZmZmZmZmZmZoiIiIiIiKqqqqqqqpmZmZmZmYiIiHd3d3d3d4iIiHd3d3d3d3d3d3d3d2ZmZlVVVURERIiIiKqqqpmZmaqqqqqqqqqqqpmZmZmZmaqqqoiIiHd3d1VVVWZmZoiIiIiIiGZmZmZmZnd3d5mZmZmZmYiIiJmZmZmZmYiIiIiIiIiIiHd3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d5mZmaqqqqqqqqqqqpmZmYiIiIiIiHd3d4iIiHd3d3d3d2ZmZnd3d3d3d3d3d0RERFVVVYiIiIiIiIiIiJmZmaqqqpmZmYiIiJmZmZmZmZmZmYiIiHd3d3d3d3d3d2ZmZmZmZlVVVWZmZoiIiHd3d3d3d5mZmYiIiIiIiIiIiHd3d4iIiHd3d3d3d3d3d3d3d2ZmZmZmZnd3d2ZmZmZmZlVVVVVVVWZmZnd3d4iIiHd3d4iIiHd3d3d3d3d3d4iIiGZmZnd3d4iIiHd3d2ZmZnd3d2ZmZmZmZmZmZlVVVVVVVURERHd3d4iIiIiIiJmZmZmZmYiIiIiIiHd3d3d3d4iIiIiIiIiIiIiIiIiIiHd3d2ZmZmZmZlVVVVVVVYiIiIiIiIiIiJmZmZmZmXd3d3d3d2ZmZmZmZlVVVVVVVWZmZlVVVWZmZlVVVWZmZmZmZmZmZlVVVURERDMzM0RERFVVVTMzMzMzM0RERFVVVTMzMyIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzM1VVVVVVVURERERERFVVVXd3d2ZmZmZmZmZmZmZmZmZmZlVVVURERFVVVVVVVVVVVURERERERERERERERERERERERFVVVURERFVVVWZmZkRERFVVVURERFVVVVVVVVVVVVVVVURERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERDMzMzMzM0RERERERERERERERGZmZnd3d1VVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVURERERERERERERERERERERERERERFVVVWZmZkRERDMzM0RERFVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzMzMzM0RERERERDMzMyIiIjMzM0RERERERERERFVVVURERFVVVURERFVVVURERFVVVURERERERERERERERDMzMzMzM0RERERERDMzM0RERDMzMzMzMzMzMyIiIkRERFVVVURERERERERERERERERERERERERERERERERERDMzM0RERDMzM0RERDMzM0RERERERERERERERERERDMzMzMzMzMzMzMzMyIiIjMzM0RERERERERERERERERERERERERERDMzM0RERDMzM0RERERERERERDMzM0RERERERERERERERERERERERERERDMzM0RERDMzMzMzMzMzMzMzMzMzM0RERFVVVURERERERERERERERERERDMzM0RERDMzM0RERERERDMzM0RERERERERERERERERERDMzM0RERFVVVVVVVVVVVVVVVVVVVURERERERERERERERERERDMzMzMzMzMzM0RERERERFVVVWZmZmZmZlVVVVVVVURERFVVVVVVVURERDMzM0RERDMzMzMzM0RERGZmZoiIiGZmZkRERFVVVXd3d2ZmZlVVVVVVVURERERERERERERERDMzM0RERFVVVURERFVVVURERERERERERERERDMzM0RERFVVVURERFVVVXd3d5mZmZmZmYiIiHd3d2ZmZlVVVVVVVVVVVVVVVURERFVVVURERERERDMzMzMzMzMzMzMzMzMzM0RERERERFVVVURERERERDMzM3d3d4iIiFVVVVVVVVVVVURERERERERERERERERERFVVVURERERERDMzMzMzMyIiIjMzMyIiIjMzMzMzM0RERDMzMyIiIjMzMzMzM0RERERERDMzMzMzMzMzM0RERERERGZmZkRERERERERERERERDMzM1VVVWZmZlVVVURERERERDMzMzMzMzMzM1VVVURERFVVVVVVVVVVVURERFVVVURERFVVVXd3d3d3d2ZmZlVVVWZmZmZmZmZmZmZmZoiIiLu7u8zMzIiIiERERDMzMyIiImZmZoiIiHd3d2ZmZlVVVURERERERDMzM0RERERERFVVVVVVVXd3d4iIiIiIiHd3d3d3d3d3d3d3d2ZmZlVVVURERERERFVVVWZmZkRERERERERERFVVVVVVVVVVVURERERERERERFVVVVVVVVVVVVVVVVVVVXd3d2ZmZlVVVVVVVVVVVWZmZmZmZnd3d5mZmYiIiIiIiIiIiHd3d5mZmZmZmWZmZjMzM0RERERERERERERERERERFVVVXd3d2ZmZlVVVVVVVWZmZnd3d0RERDMzMzMzM0RERERERERERERERFVVVWZmZmZmZmZmZmZmZkRERERERGZmZlVVVURERERERERERDMzM0RERERERERERFVVVVVVVVVVVYiIiGZmZkRERERERGZmZnd3d2ZmZmZmZlVVVVVVVVVVVVVVVURERERERERERGZmZoiIiIiIiFVVVWZmZnd3d3d3d2ZmZlVVVVVVVVVVVURERFVVVXd3d5mZmaqqqqqqqpmZmYiIiIiIiHd3d1VVVURERGZmZnd3d1VVVTMzM1VVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVXd3d5mZmXd3d3d3d3d3d5mZmXd3d2ZmZmZmZmZmZnd3d5mZmZmZmZmZmYiIiIiIiKqqqru7u7u7u6qqqru7u6qqqru7u93d3e7u7v///////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7u7u7u7u7////u7u7////u7u7////u7u7u7u7d3d3d3d3MzMzMzMzMzMzMzMy7u7vMzMy7u7vMzMy7u7uZmZmqqqqqqqrMzMzMzMzd3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3MzMzd3d3MzMzMzMzMzMzMzMzMzMy7u7u7u7uqqqqqqqqqqqqqqqqqqqqZmZmZmZmqqqqZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmIiIiZmZmIiIiIiIiZmZmIiIh3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVmZmZVVVVVVVVVVVVERERERERVVVVEREREREREREREREQzMzNEREREREREREREREQzMzMzMzMzMzMzMzNEREQzMzNERERERERERERERERERERERERVVVVERERERERVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERVVVVEREQzMzMzMzNEREQzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNEREREREQzMzMzMzNERERVVVVVVVVVVVVmZmZmZmZ3d3d3d3dmZmZVVVVVVVVmZmaIiIiIiIhVVVVVVVVERERERERmZmZmZmZ3d3eIiIiIiIh3d3dmZmZ3d3eIiIiZmZl3d3d3d3d3d3eIiIiqqqp3d3dmZmZmZmZmZmaIiIiIiIiIiIh3d3dVVVVVVVVmZmZ3d3dVVVVVVVVmZmaIiIiqqqqqqqq7u7vMzMy7u7uqqqqZmZm7u7uqqqq7u7uqqqqqqqp3d3d3d3d3d3d3d3d3d3eIiIiIiIh3d3dmZmZ3d3eZmZmZmZl3d3dVVVVmZmaqqqq7u7uIiIhmZmZmZmZ3d3d3d3dmZmZmZmZmZmZmZmZmZmaIiIh3d3d3d3d3d3eIiIiZmZmIiIiIiIiqqqqqqqqqqqqIiIiIiIiIiIh3d3eIiIiIiIh3d3d3d3dmZmZ3d3eqqqqqqqqqqqqZmZl3d3eqqqru7u7MzMy7u7u7u7uZmZmIiIiZmZmIiIiZmZmIiIh3d3eIiIiIiIiZmZmqqqqZmZmIiIiIiIiqqqrMzMyqqqqqqqqqqqqqqqq7u7uqqqqZmZmIiIiIiIh3d3eIiIiIiIiIiIiIiIhmZmZmZmZ3d3eZmZmZmZm7u7uqqqqZmZmIiIiIiIiIiIiZmZmIiIh3d3d3d3d3d3eIiIh3d3dERERmZmaqqqqZmZmIiIiZmZmqqqqZmZmZmZmZmZmIiIiIiIh3d3dmZmZ3d3eIiIh3d3dmZmZVVVVmZmaIiIiIiIh3d3eZmZmIiIiIiIh3d3eIiIh3d3dmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZ3d3eZmZmZmZmqqqqZmZmIiIiIiIiIiIiIiIh3d3d3d3dmZmZmZmZ3d3d3d3dmZmZERERVVVV3d3d3d3eIiIiZmZmIiIiZmZmIiIiZmZmIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3dVVVVmZmZ3d3dmZmaIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3dmZmZ3d3dmZmZ3d3d3d3dmZmZVVVVERERERERmZmZ3d3d3d3d3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3dmZmZmZmZmZmZmZmZVVVVERERERERmZmaIiIiIiIiIiIiIiIh3d3d3d3eIiIiIiIh3d3dmZmZ3d3eIiIiIiIh3d3dmZmZmZmZmZmZVVVVmZmZ3d3eIiIiIiIiIiIh3d3dmZmZ3d3dmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVEREREREREREREREREREQzMzNERERVVVUzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiJERERmZmZmZmYzMzMzMzNmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZERERERERERERVVVVERERVVVVVVVVVVVVVVVVVVVVERERVVVVmZmZmZmZVVVVERERVVVVERERERERVVVVmZmZVVVVERERVVVVERERVVVVVVVVVVVVVVVVERERVVVVERERVVVVEREQzMzNERERERERERERERERVVVVERERmZmZVVVVERERERERVVVVVVVVVVVVVVVVERERVVVVmZmZVVVVVVVVEREREREREREREREQzMzMzMzNVVVUzMzNERERVVVVmZmZmZmYzMzMzMzNEREQzMzNEREREREREREREREREREREREQzMzMzMzNEREQzMzNEREQzMzMzMzNERERERERERERERERERERmZmZVVVVVVVVERERVVVVEREREREREREQzMzMzMzNEREREREREREREREREREQzMzNEREQzMzMzMzNERERERERERERVVVVVVVVVVVVEREREREREREREREREREREREREREREREREREQzMzNEREQzMzNEREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNVVVVEREREREREREREREQzMzMzMzMzMzNERERERERERERERERERERVVVVEREREREREREREREQzMzMzMzNEREQzMzMzMzMzMzNEREREREREREREREREREQzMzMzMzMzMzNEREQzMzNEREQzMzNEREREREREREQzMzNEREREREREREQzMzNERERERERVVVVVVVVVVVVERERERERERERERERERERERERERERERERERERERERERERERER3d3dmZmYzMzNERERVVVVVVVVEREREREREREQzMzMzMzMzMzMzMzN3d3eqqqp3d3dVVVVVVVVVVVVmZmZVVVVEREREREREREREREQzMzMzMzNERERVVVVmZmZVVVVVVVVEREREREQzMzNERERmZmZmZmZERERVVVVmZmaZmZmZmZl3d3dmZmZmZmZVVVVERERVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERERERVVVV3d3dmZmZVVVVVVVV3d3dmZmZVVVVERERERERERERERERVVVVVVVVEREQzMzMzMzMzMzMiIiIzMzMzMzNEREQzMzMzMzMzMzMzMzNEREREREQzMzMiIiIzMzMzMzNERERVVVVEREREREREREQzMzNERERVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERERERVVVVERERERERERERERERVVVV3d3d3d3dmZmZVVVVmZmZmZmZmZmZmZmaIiIjMzMzMzMx3d3dEREQzMzMiIiJVVVV3d3d3d3d3d3dmZmZEREREREREREQzMzNERERERERmZmaIiIh3d3eIiIh3d3d3d3d3d3eIiIiZmZlmZmZVVVVVVVVmZmZVVVVEREQzMzMzMzNVVVVERERERERERERVVVVERERVVVVVVVVVVVVVVVVVVVV3d3eIiIhVVVVVVVVERERVVVV3d3dmZmZ3d3d3d3dmZmZmZmZ3d3eIiIiZmZlmZmZEREREREQzMzNERERmZmZVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZVVVVERERERERVVVVVVVVERERERERVVVVmZmZmZmZVVVVEREQzMzMzMzNEREREREREREQzMzMzMzNERERERERVVVVVVVVmZmZmZmaIiIiqqqp3d3dERERERERmZmZmZmZmZmZmZmZmZmZVVVVVVVVERERERERERERVVVVVVVVmZmZmZmZVVVVmZmaIiIh3d3d3d3dVVVVmZmZmZmZVVVVERERVVVVmZmZ3d3eIiIhmZmZVVVVEREREREQzMzNERERVVVVVVVUzMzNERER3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZ3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3dmZmZVVVVVVVVVVVVmZmaZmZmqqqqZmZmZmZmIiIiZmZmqqqqZmZmqqqqqqqrMzMy7u7vMzMz///////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u////7u7u////7u7u7u7u7u7u////7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u7u7u3d3d7u7u3d3d7u7u3d3d3d3d3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzMzMzMzMzMzMzMu7u7qqqqqqqqqqqqmZmZiIiImZmZiIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3ZmZmd3d3d3d3ZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmVVVVREREREREREREVVVVREREVVVVREREREREREREREREREREREREREREREREREREREREREREREREMzMzMzMzREREREREREREMzMzREREREREMzMzREREREREMzMzMzMzMzMzREREREREREREREREREREMzMzREREREREREREREREREREREREREREREREREREVVVVREREREREREREVVVVREREMzMzMzMzREREREREREREMzMzREREMzMzMzMzVVVVVVVVREREVVVVREREREREREREVVVVREREREREREREVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmVVVVZmZmZmZmZmZmZmZmd3d3ZmZmZmZmVVVVVVVVVVVVd3d3ZmZmVVVVREREREREVVVVVVVVZmZmd3d3d3d3d3d3ZmZmiIiImZmZiIiId3d3d3d3iIiIqqqqmZmZd3d3ZmZmZmZmiIiIiIiIiIiId3d3ZmZmVVVVZmZmZmZmd3d3ZmZmVVVVZmZmmZmZqqqqzMzMzMzMzMzMqqqqqqqqqqqqu7u7zMzMu7u7qqqqqqqqiIiIiIiIiIiId3d3d3d3d3d3iIiImZmZiIiId3d3iIiImZmZd3d3ZmZmd3d3mZmZmZmZmZmZd3d3d3d3d3d3ZmZmd3d3ZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3iIiImZmZiIiImZmZmZmZiIiIiIiIiIiIiIiIiIiId3d3d3d3iIiIiIiId3d3d3d3iIiImZmZqqqqqqqqiIiIiIiIzMzM3d3dzMzMu7u7qqqqmZmZiIiId3d3iIiId3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIqqqqu7u7u7u7mZmZqqqqqqqqqqqqqqqqqqqqqqqqmZmZd3d3iIiIiIiIiIiImZmZiIiIZmZmVVVViIiImZmZqqqqqqqqmZmZiIiIqqqqmZmZmZmZiIiIiIiIiIiId3d3iIiId3d3ZmZmVVVVd3d3mZmZmZmZiIiId3d3iIiImZmZiIiImZmZiIiIiIiId3d3ZmZmd3d3d3d3ZmZmZmZmVVVVZmZmiIiId3d3d3d3mZmZmZmZiIiIiIiIiIiId3d3ZmZmVVVVZmZmZmZmZmZmd3d3ZmZmVVVVZmZmiIiImZmZmZmZiIiImZmZiIiIiIiIiIiId3d3ZmZmd3d3ZmZmd3d3ZmZmZmZmREREREREZmZmd3d3iIiIiIiId3d3iIiId3d3iIiIiIiIiIiIiIiId3d3iIiId3d3d3d3ZmZmVVVVVVVVd3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3ZmZmREREREREZmZmd3d3d3d3ZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmVVVVZmZmREREREREREREZmZmiIiId3d3d3d3d3d3iIiId3d3d3d3iIiId3d3ZmZmd3d3d3d3iIiId3d3ZmZmZmZmZmZmVVVVVVVVZmZmiIiIiIiIiIiId3d3ZmZmZmZmd3d3ZmZmZmZmZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREREREMzMzREREMzMzREREREREREREMzMzIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzVVVVVVVVMzMzREREVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREZmZmd3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmZmZmREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREREREMzMzREREVVVVREREREREVVVVVVVVREREVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREMzMzMzMzMzMzREREMzMzREREREREZmZmVVVVVVVVREREREREMzMzREREREREREREMzMzREREREREREREMzMzMzMzMzMzREREMzMzIiIiREREVVVVREREREREREREVVVVVVVVREREVVVVREREREREREREMzMzREREREREREREREREREREREREVVVVREREMzMzMzMzMzMzVVVVREREREREREREVVVVVVVVVVVVREREREREREREREREMzMzREREMzMzMzMzREREREREREREREREREREREREREREREREMzMzREREMzMzMzMzMzMzREREREREREREREREREREREREREREREREMzMzMzMzREREREREREREREREREREREREVVVVREREREREREREREREMzMzMzMzMzMzMzMzMzMzREREVVVVREREREREMzMzMzMzREREMzMzREREMzMzREREREREREREREREREREREREREREREREMzMzMzMzMzMzVVVVVVVVZmZmVVVVREREREREMzMzREREREREREREREREMzMzREREREREMzMzREREVVVVVVVVREREREREVVVVVVVVREREMzMzREREMzMzIiIiMzMzMzMzVVVViIiIiIiIZmZmVVVVZmZmVVVVREREZmZmVVVVVVVVREREREREREREREREVVVVVVVVVVVVREREVVVVREREMzMzREREd3d3VVVVREREVVVVZmZmiIiIqqqqd3d3d3d3d3d3VVVVREREVVVVVVVVMzMzREREMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVd3d3VVVVREREVVVVd3d3d3d3VVVVVVVVVVVVREREREREREREREREVVVVREREMzMzMzMzIiIiMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzREREMzMzMzMzREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREMzMzREREREREREREREREMzMzREREVVVVZmZmiIiIiIiIZmZmZmZmZmZmZmZmd3d3ZmZmmZmZzMzMzMzMd3d3REREMzMzIiIiVVVVd3d3ZmZmZmZmVVVVVVVVVVVVREREMzMzREREVVVVd3d3d3d3d3d3iIiIiIiIZmZmd3d3mZmZmZmZZmZmd3d3ZmZmZmZmVVVVMzMzMzMzREREREREREREREREREREVVVVREREREREVVVVVVVVVVVVZmZmZmZmd3d3VVVVVVVVVVVVVVVVZmZmZmZmVVVVZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmREREREREREREREREVVVVREREVVVVVVVVZmZmiIiId3d3VVVVVVVVREREREREVVVVVVVVREREVVVVZmZmZmZmVVVVVVVVREREREREMzMzMzMzREREVVVVREREREREREREVVVVZmZmZmZmZmZmmZmZqqqqzMzMiIiIREREVVVVZmZmZmZmZmZmd3d3ZmZmVVVVREREREREVVVVVVVVREREREREVVVVVVVVVVVVVVVVd3d3d3d3d3d3ZmZmd3d3d3d3VVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREMzMzVVVVZmZmZmZmMzMzIiIiVVVVd3d3iIiIiIiIiIiIiIiIiIiImZmZmZmZmZmZqqqqqqqqmZmZmZmZmZmZiIiImZmZmZmZiIiId3d3d3d3d3d3ZmZmVVVVZmZmZmZmd3d3d3d3iIiIiIiIiIiIiIiImZmZmZmZmZmZmZmZqqqqzMzMzMzM3d3d////7u7u////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3e7u7t3d3e7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3d3d3d3d3e7u7t3d3e7u7t3d3d3d3d3d3czMzMzMzLu7u7u7u6qqqqqqqpmZmZmZmXd3d3d3d2ZmZlVVVWZmZmZmZlVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERERERERERERERERERERERERERERERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERDMzMzMzM0RERDMzMzMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERDMzMzMzM0RERGZmZmZmZlVVVVVVVVVVVURERFVVVWZmZmZmZlVVVVVVVWZmZlVVVWZmZnd3d3d3d1VVVVVVVXd3d1VVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVWZmZnd3d2ZmZmZmZlVVVWZmZmZmZlVVVXd3d3d3d2ZmZnd3d2ZmZnd3d4iIiHd3d3d3d6qqqqqqqnd3d2ZmZoiIiIiIiIiIiIiIiIiIiIiIiHd3d2ZmZmZmZmZmZnd3d2ZmZmZmZpmZmZmZmaqqqszMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u6qqqpmZmYiIiJmZmYiIiJmZmZmZmYiIiHd3d4iIiJmZmYiIiGZmZnd3d3d3d3d3d4iIiJmZmZmZmYiIiJmZmYiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d3d3d3d3d5mZmYiIiJmZmZmZmYiIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiIiIiIiIiIiIiJmZmZmZmZmZmYiIiIiIiKqqqszMzMzMzLu7u6qqqqqqqpmZmYiIiIiIiIiIiHd3d4iIiHd3d4iIiJmZmXd3d2ZmZnd3d4iIiJmZmaqqqru7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqpmZmYiIiIiIiJmZmYiIiHd3d3d3d1VVVWZmZpmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmYiIiHd3d3d3d3d3d2ZmZmZmZmZmZlVVVXd3d4iIiJmZmYiIiIiIiJmZmZmZmYiIiIiIiIiIiHd3d3d3d3d3d3d3d2ZmZmZmZmZmZkRERGZmZnd3d3d3d5mZmZmZmYiIiIiIiHd3d3d3d3d3d2ZmZnd3d2ZmZmZmZnd3d3d3d2ZmZlVVVWZmZoiIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiHd3d2ZmZnd3d3d3d2ZmZlVVVVVVVURERERERGZmZnd3d4iIiIiIiIiIiHd3d3d3d4iIiHd3d3d3d3d3d4iIiHd3d3d3d2ZmZnd3d1VVVWZmZnd3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZnd3d3d3d3d3d2ZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZlVVVURERERERERERGZmZnd3d2ZmZnd3d4iIiHd3d4iIiIiIiIiIiHd3d2ZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVWZmZmZmZnd3d4iIiHd3d2ZmZlVVVWZmZnd3d3d3d2ZmZlVVVVVVVVVVVVVVVWZmZlVVVVVVVURERERERDMzM0RERDMzMzMzM0RERERERDMzMyIiIjMzMzMzM0RERERERERERDMzMzMzMzMzM0RERDMzM0RERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVXd3d2ZmZmZmZnd3d3d3d3d3d2ZmZlVVVWZmZnd3d3d3d1VVVWZmZlVVVURERERERERERFVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVURERFVVVURERERERERERERERERERFVVVURERERERFVVVURERERERFVVVURERERERERERERERDMzM0RERERERERERERERERERERERERERERERFVVVURERFVVVVVVVVVVVURERERERDMzMzMzMzMzMzMzM0RERDMzM0RERERERERERCIiIjMzMzMzM0RERERERDMzM0RERERERERERDMzM0RERERERERERERERDMzM0RERERERFVVVVVVVURERFVVVURERERERERERDMzM0RERERERERERERERERERFVVVURERFVVVURERERERERERERERDMzM0RERERERERERERERERERERERFVVVVVVVURERERERDMzM0RERDMzMzMzMzMzMzMzMzMzM0RERFVVVURERERERERERDMzMzMzM0RERDMzMzMzM0RERDMzM0RERERERERERERERDMzM0RERDMzM0RERDMzMzMzMzMzMzMzMzMzM0RERERERFVVVURERERERERERERERERERDMzM0RERERERERERERERERERERERDMzM0RERERERDMzMzMzMzMzM2ZmZmZmZmZmZlVVVURERDMzMzMzM0RERERERERERERERERERDMzM0RERDMzMzMzM0RERERERERERERERFVVVWZmZkRERDMzMzMzMzMzMzMzMzMzMzMzMzMzM2ZmZnd3d1VVVWZmZnd3d1VVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERDMzM2ZmZnd3d1VVVVVVVVVVVVVVVXd3d4iIiIiIiHd3d2ZmZlVVVVVVVURERERERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERGZmZnd3d1VVVURERGZmZnd3d3d3d1VVVVVVVVVVVURERERERDMzM0RERERERERERDMzMyIiIjMzMzMzMzMzM0RERERERDMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzM1VVVVVVVVVVVWZmZlVVVVVVVURERFVVVVVVVURERERERERERERERERERDMzM0RERERERFVVVXd3d4iIiIiIiGZmZmZmZmZmZnd3d3d3d2ZmZpmZmczMzMzMzHd3d0RERERERCIiIlVVVYiIiHd3d2ZmZlVVVURERFVVVVVVVURERFVVVWZmZnd3d2ZmZnd3d3d3d4iIiHd3d4iIiJmZmYiIiGZmZmZmZmZmZlVVVVVVVTMzMzMzMzMzMzMzM0RERERERERERERERERERFVVVVVVVVVVVWZmZlVVVVVVVWZmZmZmZkRERFVVVWZmZlVVVVVVVVVVVVVVVWZmZlVVVVVVVWZmZmZmZnd3d2ZmZlVVVURERERERERERERERERERFVVVVVVVWZmZoiIiHd3d2ZmZmZmZkRERERERERERERERFVVVVVVVVVVVVVVVWZmZmZmZmZmZkRERERERERERFVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZoiIiJmZmbu7u3d3d0RERFVVVWZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVURERFVVVURERFVVVVVVVWZmZmZmZnd3d2ZmZlVVVVVVVXd3d3d3d0RERERERERERERERDMzM0RERGZmZoiIiGZmZjMzMzMzM3d3d4iIiIiIiIiIiIiIiIiIiJmZmZmZmaqqqru7u8zMzO7u7szMzN3d3czMzMzMzMzMzMzMzLu7u6qqqpmZmYiIiJmZmYiIiGZmZmZmZmZmZmZmZoiIiIiIiIiIiIiIiKqqqpmZmaqqqqqqqru7u8zMzO7u7v///////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////u7u7d3d3d3d3d3d3d3d3MzMzMzMzd3d3MzMzMzMzMzMzMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7d3d3d3d3u7u7d3d3d3d3d3d3MzMzMzMy7u7u7u7uqqqqZmZmIiIiIiIh3d3dmZmZmZmZVVVVVVVVEREREREREREQzMzNEREQzMzNEREQzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIzMzMiIiIiIiIiIiIzMzNEREQzMzMzMzNEREREREQzMzMzMzNEREQzMzNEREQzMzMiIiIzMzMzMzMzMzMzMzNEREREREREREQzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzNERERERERERERmZmZVVVVERERERERVVVVERERERERERERERERVVVVVVVV3d3dmZmZERERERERVVVVERERERERERERVVVVERERVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3eIiIh3d3dVVVVmZmZ3d3eIiIiIiIh3d3dmZmZmZmZ3d3eIiIiqqqqZmZlmZmaIiIiZmZmZmZmZmZmZmZmIiIh3d3eIiIiIiIiIiIiIiIh3d3dERERmZmaZmZnMzMzMzMy7u7u7u7u7u7vMzMy7u7u7u7u7u7u7u7uZmZmIiIiIiIiZmZmZmZmqqqqqqqqZmZmZmZmIiIiZmZmIiIiIiIh3d3dmZmaIiIiZmZmZmZmZmZmZmZmIiIiZmZmIiIiIiIiIiIiIiIh3d3d3d3eIiIh3d3d3d3d3d3d3d3dmZmZmZmaZmZmqqqq7u7uqqqqqqqqqqqqZmZmIiIiIiIiZmZmIiIiIiIiIiIiZmZmZmZmZmZmZmZmIiIh3d3eIiIi7u7vMzMzMzMyqqqqqqqqqqqqZmZmIiIiIiIiIiIiZmZl3d3d3d3eIiIiIiIhmZmZmZmZ3d3d3d3eIiIiZmZm7u7u7u7uZmZmqqqqqqqqqqqqqqqqZmZmZmZmZmZmIiIiIiIiIiIhmZmZVVVVmZmZmZmaIiIiZmZmZmZmZmZmZmZmZmZmIiIh3d3eIiIiIiIhmZmZmZmZVVVVVVVVmZmZ3d3dVVVV3d3eIiIiIiIiZmZmZmZmZmZmZmZmIiIiIiIiIiIh3d3dmZmZ3d3dmZmZmZmZ3d3dVVVVVVVVERER3d3d3d3eIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZVVVVVVVVmZmZ3d3eIiIiIiIh3d3d3d3d3d3d3d3dmZmZmZmZmZmZ3d3d3d3dmZmZVVVVVVVVVVVVERERmZmaIiIh3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3eIiIiIiIh3d3d3d3d3d3dmZmZVVVV3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZ3d3d3d3dmZmZmZmZ3d3d3d3d3d3dmZmZmZmZ3d3dmZmZVVVVVVVVmZmZmZmZVVVVVVVVERERVVVVmZmZmZmZVVVVVVVVVVVVVVVVmZmZVVVVmZmZVVVVVVVVERERERERERERmZmZVVVVmZmZ3d3d3d3d3d3eIiIiIiIiIiIh3d3d3d3d3d3d3d3dmZmZ3d3dmZmZ3d3dmZmZERERERERVVVVmZmZ3d3d3d3dVVVVVVVVmZmZVVVVmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVEREREREQzMzMzMzMzMzMzMzNEREREREREREQzMzMiIiIzMzNERERVVVVERERERERERERERERERERERERVVVVmZmZ3d3dmZmZ3d3dmZmZmZmZVVVV3d3dmZmZVVVVERERVVVVVVVVERERVVVVmZmZmZmZVVVVVVVV3d3eIiIiIiIh3d3eIiIh3d3dmZmaIiIh3d3d3d3eIiIiIiIhVVVVVVVVVVVVVVVVERERERERmZmZ3d3dmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZVVVVmZmZVVVVVVVVVVVVVVVVEREREREREREREREQzMzNEREQzMzNEREQzMzNERERERERVVVVERERERERVVVVERERVVVVVVVVVVVVERERERERERERVVVVVVVVVVVVEREREREREREQzMzMzMzMzMzNERERVVVVEREREREQzMzMzMzNEREREREREREREREREREREREREREQzMzNEREQzMzMzMzNERERERERVVVVVVVVVVVVERERVVVVEREREREREREREREREREREREREREREREQzMzNERERERERVVVVERERERERERERERERERERERERERERERERERERERERERERVVVVERERVVVVEREREREREREREREREREQzMzNEREQzMzMzMzNEREREREREREREREREREREREQzMzNEREQzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMiIiIiIiIzMzNERERERERERERVVVVVVVVEREREREQzMzNEREREREQzMzNEREREREREREREREREREREREQzMzNEREQzMzNERERVVVVVVVVVVVVVVVVVVVVEREREREQzMzNEREREREREREREREREREREREQzMzMzMzNERERVVVVVVVVERERVVVVVVVUzMzNEREQzMzNEREQzMzMzMzNERERVVVWIiIhmZmZmZmZmZmaIiIiIiIhmZmZVVVVVVVVVVVVERERERERERERVVVVERERVVVVEREREREREREREREQzMzNVVVVmZmZERERERERERERVVVVmZmaIiIiIiIhmZmZmZmZVVVVERERERERERERERERVVVVERERVVVVEREREREQzMzMzMzMiIiIzMzMzMzMzMzMzMzNERERmZmZmZmZVVVVVVVVmZmZ3d3dVVVVVVVVmZmZVVVVEREQzMzNEREREREREREQzMzMiIiIzMzMzMzMzMzMzMzMzMzNEREQzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIzMzMiIiIzMzNERERVVVVERERERERVVVVVVVVERERERERVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVV3d3eIiIiIiIh3d3eIiIiIiIh3d3eIiIh3d3eIiIi7u7vMzMx3d3dVVVVEREQzMzNERESIiIiZmZmIiIhmZmZERERVVVVVVVVVVVVVVVVVVVVERERERERVVVVmZmZ3d3eIiIiZmZmIiIh3d3dmZmZVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzNERERERERERERVVVVERERVVVVVVVVVVVVmZmZ3d3dmZmZmZmZmZmZVVVVERERERERVVVVVVVVVVVVmZmZmZmZmZmZERERERERmZmZmZmZmZmZmZmZVVVVERERERERVVVVVVVVERERmZmZmZmZVVVV3d3eIiIhmZmZVVVVVVVVERERERERVVVVVVVVERERERERVVVVmZmZmZmZVVVV3d3dmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3d3d3d3d3eIiIhmZmZVVVVERERVVVVmZmZ3d3dmZmZVVVVVVVVVVVVVVVWIiIiqqqp3d3dVVVVVVVVVVVVERERVVVVERERERERERERVVVVVVVVVVVVmZmZVVVVmZmZmZmZEREQzMzMzMzNERERERERVVVV3d3eIiIhVVVUzMzNVVVVmZmaIiIiIiIh3d3eIiIiIiIiIiIiIiIiqqqrd3d3d3d3u7u7u7u7u7u7u7u7u7u7d3d3d3d3MzMzMzMzMzMy7u7u7u7u7u7uZmZmIiIiIiIh3d3d3d3eIiIiIiIiZmZmZmZmZmZmqqqq7u7vMzMzu7u7////u7u7u7u7///////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u3d3d3d3d3d3d3d3dzMzM3d3dzMzM3d3d3d3d3d3d3d3d7u7u3d3d7u7u3d3d7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3dzMzMzMzMzMzMzMzM3d3dzMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7qqqqqqqqqqqqmZmZmZmZiIiIiIiId3d3d3d3d3d3d3d3ZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiMzMzMzMzMzMzIiIiMzMzREREMzMzMzMzREREREREMzMzREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzMzMzREREMzMzMzMzMzMzREREMzMzREREVVVVVVVVREREREREVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmVVVVZmZmZmZmZmZmZmZmd3d3d3d3iIiIiIiIiIiIZmZmZmZmiIiImZmZiIiIiIiId3d3ZmZmZmZmd3d3mZmZmZmZd3d3iIiIiIiIiIiIiIiImZmZiIiId3d3iIiIiIiIiIiId3d3d3d3VVVViIiIqqqqzMzMzMzMzMzMqqqqqqqqqqqqqqqqqqqqzMzMqqqqmZmZmZmZmZmZmZmZqqqqqqqqqqqqqqqqmZmZmZmZiIiIiIiId3d3ZmZmZmZmiIiImZmZiIiImZmZiIiImZmZiIiIiIiIiIiIiIiIiIiImZmZiIiIiIiIiIiId3d3d3d3d3d3ZmZmZmZmmZmZqqqqqqqqqqqqqqqqqqqqqqqqiIiImZmZiIiImZmZmZmZmZmZmZmZmZmZiIiIiIiId3d3ZmZmmZmZu7u7zMzMu7u7qqqqiIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3iIiIiIiId3d3d3d3ZmZmiIiId3d3iIiIqqqqu7u7qqqqqqqqqqqqqqqqmZmZmZmZmZmZiIiIiIiIiIiIiIiId3d3ZmZmREREVVVVd3d3iIiIqqqqmZmZqqqqqqqqiIiIiIiId3d3d3d3iIiId3d3VVVVZmZmZmZmVVVVVVVVVVVVd3d3mZmZmZmZiIiIiIiId3d3iIiId3d3iIiId3d3ZmZmd3d3d3d3ZmZmZmZmVVVVVVVVREREVVVVd3d3d3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmVVVVVVVVZmZmZmZmd3d3iIiId3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmd3d3ZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmd3d3d3d3d3d3iIiIiIiId3d3d3d3d3d3ZmZmZmZmVVVVd3d3ZmZmd3d3ZmZmZmZmd3d3ZmZmd3d3d3d3d3d3ZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVMzMzMzMzREREVVVVVVVVZmZmd3d3d3d3d3d3iIiIiIiId3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3ZmZmVVVVREREVVVVd3d3d3d3ZmZmZmZmd3d3d3d3d3d3ZmZmVVVVZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmREREREREVVVVREREREREREREZmZmVVVVREREMzMzMzMzMzMzREREVVVVREREVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVZmZmZmZmVVVVZmZmd3d3ZmZmZmZmVVVVVVVVREREVVVVREREVVVVVVVVVVVVREREZmZmZmZmZmZmd3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVREREREREREREREREVVVVREREREREREREREREREREREREREREREREVVVVREREREREREREVVVVREREREREVVVVVVVVVVVVREREREREMzMzIiIiREREVVVVREREREREREREMzMzREREREREREREREREREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREMzMzREREVVVVVVVVREREREREREREMzMzREREMzMzREREREREMzMzREREREREREREREREVVVVVVVVREREVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzREREREREREREREREREREREREMzMzREREREREREREREREREREREREREREMzMzMzMzREREREREMzMzREREREREREREREREREREREREREREREREREREREREREREREREREREREREMzMzMzMzREREREREZmZmVVVVVVVVREREREREREREMzMzMzMzREREMzMzMzMzREREiIiImZmZZmZmZmZmZmZmd3d3iIiId3d3ZmZmVVVVREREREREREREREREREREREREVVVVREREVVVVVVVVREREMzMzREREREREMzMzMzMzREREVVVVZmZmmZmZmZmZd3d3ZmZmVVVVREREVVVVVVVVREREREREREREVVVVVVVVVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzVVVVZmZmVVVVZmZmZmZmd3d3ZmZmVVVVVVVVZmZmVVVVREREMzMzMzMzREREREREMzMzMzMzMzMzMzMzREREREREREREREREMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzREREREREMzMzREREVVVVREREVVVVVVVVVVVVREREREREREREVVVVVVVVZmZmZmZmZmZmd3d3ZmZmZmZmd3d3iIiIiIiIiIiId3d3iIiImZmZd3d3d3d3qqqqu7u7iIiIVVVVMzMzIiIiREREmZmZqqqqiIiIZmZmZmZmVVVVVVVVREREREREREREMzMzREREREREVVVViIiImZmZmZmZmZmZmZmZd3d3ZmZmVVVVVVVVREREMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVVVVVVVVVVVVVd3d3d3d3d3d3VVVVZmZmVVVVREREREREREREVVVVZmZmZmZmVVVVVVVVREREREREZmZmVVVVZmZmVVVVVVVVREREVVVVREREREREVVVVVVVVVVVVZmZmZmZmiIiId3d3ZmZmVVVVREREREREVVVVREREREREREREREREVVVVZmZmZmZmiIiId3d3ZmZmVVVVVVVVZmZmZmZmVVVVZmZmd3d3ZmZmZmZmZmZmd3d3ZmZmREREVVVVVVVVd3d3iIiId3d3VVVVVVVVVVVVVVVVd3d3mZmZd3d3VVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3ZmZmVVVVREREREREREREVVVVVVVVZmZmZmZmd3d3REREREREVVVVZmZmd3d3d3d3d3d3iIiIiIiIiIiIiIiIu7u73d3d3d3d7u7u3d3d3d3d7u7u3d3d3d3dzMzMu7u7zMzMu7u7qqqqqqqqqqqqu7u7qqqqqqqqqqqqmZmZmZmZmZmZmZmZmZmZmZmZqqqq3d3d3d3d3d3d7u7uzMzM3d3d////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////+7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7u7u7t3d3d3d3czMzLu7u6qqqpmZmZmZmZmZmaqqqqqqqqqqqqqqqqqqqqqqqru7u7u7u7u7u7u7u7u7u7u7u6qqqpmZmaqqqpmZmaqqqpmZmZmZmZmZmYiIiHd3d2ZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZlVVVVVVVWZmZlVVVVVVVVVVVVVVVURERFVVVVVVVURERERERFVVVURERERERERERERERERERERERFVVVURERERERERERERERDMzM0RERERERERERFVVVURERERERERERERERERERDMzM0RERDMzMzMzMzMzM0RERDMzM0RERDMzM0RERDMzM0RERERERERERERERERERERERFVVVVVVVVVVVURERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM0RERDMzMzMzM0RERERERFVVVURERFVVVURERERERFVVVWZmZnd3d2ZmZlVVVVVVVVVVVWZmZmZmZlVVVWZmZlVVVVVVVXd3d3d3d3d3d4iIiIiIiHd3d4iIiIiIiHd3d4iIiJmZmYiIiJmZmZmZmWZmZnd3d4iIiIiIiIiIiHd3d4iIiIiIiHd3d3d3d4iIiIiIiHd3d2ZmZmZmZoiIiHd3d2ZmZnd3d7u7u8zMzMzMzMzMzLu7u7u7u5mZmYiIiJmZmbu7u7u7u5mZmZmZmaqqqpmZmaqqqpmZmaqqqqqqqqqqqpmZmYiIiIiIiIiIiGZmZlVVVWZmZoiIiIiIiJmZmYiIiJmZmYiIiHd3d4iIiHd3d4iIiIiIiHd3d4iIiIiIiIiIiIiIiHd3d4iIiGZmZmZmZqqqqqqqqpmZmYiIiKqqqpmZmaqqqpmZmYiIiIiIiJmZmZmZmZmZmYiIiJmZmZmZmYiIiGZmZmZmZpmZmbu7u7u7u6qqqoiIiHd3d4iIiHd3d3d3d3d3d2ZmZmZmZnd3d3d3d3d3d3d3d3d3d4iIiIiIiGZmZoiIiKqqqru7u6qqqqqqqpmZmYiIiJmZmYiIiIiIiHd3d3d3d4iIiHd3d4iIiGZmZlVVVVVVVXd3d4iIiJmZmaqqqpmZmZmZmYiIiIiIiHd3d4iIiHd3d4iIiHd3d2ZmZlVVVVVVVURERFVVVWZmZpmZmZmZmZmZmYiIiHd3d3d3d3d3d4iIiGZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVURERFVVVXd3d4iIiIiIiHd3d2ZmZmZmZnd3d3d3d3d3d3d3d3d3d2ZmZlVVVVVVVWZmZmZmZnd3d3d3d3d3d4iIiHd3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZlVVVVVVVVVVVURERFVVVVVVVXd3d1VVVWZmZmZmZnd3d2ZmZnd3d3d3d4iIiIiIiIiIiIiIiHd3d3d3d2ZmZmZmZmZmZmZmZnd3d3d3d3d3d1VVVVVVVWZmZnd3d2ZmZnd3d2ZmZmZmZnd3d3d3d2ZmZmZmZmZmZlVVVVVVVURERERERGZmZnd3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d2ZmZmZmZlVVVURERERERDMzM0RERDMzM1VVVWZmZoiIiIiIiHd3d3d3d4iIiHd3d3d3d2ZmZmZmZnd3d2ZmZmZmZnd3d3d3d2ZmZkRERERERFVVVWZmZnd3d3d3d3d3d2ZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZpmZmZmZmYiIiIiIiHd3d2ZmZnd3d2ZmZlVVVURERFVVVVVVVVVVVVVVVURERERERERERFVVVURERFVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVURERFVVVVVVVVVVVVVVVXd3d3d3d4iIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d3d3d2ZmZnd3d3d3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVWZmZlVVVVVVVURERERERFVVVWZmZlVVVURERERERERERERERFVVVURERDMzM0RERGZmZlVVVURERERERDMzMzMzMzMzM0RERFVVVURERERERERERERERERERERERERERERERERERERERDMzM0RERERERERERERERERERERERFVVVURERERERERERERERERERERERERERFVVVURERDMzM0RERERERFVVVVVVVURERERERERERERERERERDMzM0RERERERERERERERERERERERDMzM0RERDMzMzMzM0RERDMzMzMzMzMzM0RERFVVVURERERERERERFVVVWZmZlVVVURERDMzM0RERDMzMzMzM0RERDMzMzMzMyIiIjMzMyIiIjMzMzMzM0RERDMzMzMzMzMzMyIiIjMzMyIiIjMzM0RERERERERERFVVVURERDMzM0RERERERDMzM0RERERERDMzM0RERERERERERERERERERERERERERDMzM0RERERERFVVVVVVVURERERERERERERERDMzM0RERDMzMzMzM0RERDMzM0RERERERFVVVWZmZlVVVURERERERERERDMzMyIiIjMzMzMzM0RERDMzM0RERIiIiIiIiFVVVVVVVWZmZnd3d3d3d4iIiFVVVURERERERERERERERFVVVURERERERERERERERFVVVURERERERDMzM0RERFVVVTMzMzMzM0RERFVVVWZmZpmZmZmZmYiIiHd3d2ZmZlVVVWZmZlVVVWZmZlVVVURERERERERERFVVVVVVVURERERERDMzM0RERDMzMzMzM1VVVWZmZmZmZnd3d3d3d3d3d2ZmZlVVVVVVVVVVVVVVVURERERERDMzM0RERERERDMzMyIiIjMzMzMzM0RERERERERERFVVVURERERERERERDMzMyIiIiIiIiIiIjMzMzMzMyIiIjMzM0RERFVVVVVVVURERERERERERERERDMzM0RERFVVVVVVVVVVVURERERERFVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVXd3d4iIiIiIiHd3d4iIiIiIiJmZmYiIiHd3d5mZmczMzJmZmVVVVURERCIiIkRERIiIiIiIiHd3d2ZmZlVVVVVVVVVVVURERERERDMzM0RERERERERERERERHd3d4iIiKqqqpmZmYiIiGZmZlVVVVVVVXd3d1VVVTMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVURERFVVVVVVVVVVVYiIiIiIiGZmZlVVVWZmZlVVVURERERERERERERERERERERERERERERERFVVVWZmZmZmZlVVVVVVVURERERERERERERERFVVVVVVVVVVVVVVVWZmZmZmZnd3d4iIiHd3d1VVVVVVVVVVVURERFVVVVVVVURERFVVVVVVVWZmZnd3d3d3d4iIiGZmZlVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVWZmZoiIiHd3d1VVVURERFVVVXd3d3d3d3d3d2ZmZlVVVVVVVXd3d3d3d3d3d3d3d2ZmZlVVVWZmZlVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVWZmZnd3d2ZmZkRERDMzM0RERGZmZnd3d2ZmZlVVVWZmZlVVVURERERERGZmZnd3d2ZmZnd3d2ZmZnd3d3d3d5mZmbu7u8zMzLu7u93d3f///93d3d3d3czMzMzMzLu7u6qqqqqqqqqqqru7u6qqqqqqqpmZmZmZmaqqqru7u6qqqru7u7u7u6qqqqqqqru7u6qqqru7u93d3d3d3d3d3czMzMzMzO7u7v///////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////u7u7////u7u7u7u7d3d3u7u7d3d3MzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7uqqqqqqqqqqqqqqqqqqqq7u7u7u7vMzMy7u7vMzMyqqqqqqqqZmZmZmZmZmZmZmZmIiIiZmZmqqqq7u7vMzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3MzMy7u7vMzMy7u7u7u7uqqqq7u7uqqqqqqqqZmZmZmZmqqqqZmZmZmZmqqqqZmZmZmZmqqqqZmZmZmZmZmZmIiIh3d3eIiIiIiIiIiIiIiIiIiIh3d3eIiIiIiIiIiIh3d3d3d3eIiIiIiIh3d3d3d3d3d3dmZmZ3d3d3d3dmZmZ3d3d3d3d3d3dmZmZ3d3dmZmZmZmZ3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZmZmZ3d3dmZmZVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZVVVVVVVVmZmZ3d3eIiIh3d3eIiIiZmZmIiIiZmZmZmZmIiIiIiIiZmZmZmZmZmZmZmZmIiIiIiIiZmZmIiIiIiIh3d3eIiIiIiIh3d3eIiIiIiIh3d3d3d3d3d3eIiIh3d3dVVVVVVVW7u7vd3d3d3d3MzMzMzMzMzMy7u7uqqqqIiIiqqqrMzMyqqqqqqqqZmZmZmZmqqqq7u7uqqqqZmZmqqqqZmZmZmZmZmZmZmZl3d3dmZmZmZmZ3d3eIiIiZmZmIiIiIiIh3d3d3d3eIiIiIiIiIiIiIiIh3d3d3d3eIiIiIiIiIiIh3d3eIiIiIiIhmZmZmZmaZmZmqqqqZmZmIiIiZmZmZmZmIiIiIiIiZmZmIiIiZmZmZmZmZmZmZmZmZmZmIiIh3d3dmZmZ3d3eZmZmqqqqZmZmIiIiIiIh3d3dmZmZ3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3eIiIiqqqqqqqqZmZmIiIiZmZmIiIh3d3d3d3eIiIh3d3eIiIh3d3d3d3d3d3dmZmZVVVVVVVVmZmaIiIiIiIiIiIiIiIiIiIh3d3dmZmZ3d3d3d3eIiIh3d3eIiIhmZmZmZmZERERVVVVVVVVVVVV3d3eZmZmIiIh3d3d3d3d3d3d3d3d3d3dmZmZVVVVmZmZmZmZVVVVVVVVVVVVERERVVVVmZmZmZmZ3d3d3d3d3d3dmZmZ3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVERERVVVVVVVVERERVVVVmZmZmZmZmZmZmZmZ3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3dVVVVmZmZ3d3dmZmZmZmZVVVVVVVVmZmZmZmZVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZVVVVEREQzMzNERERmZmZmZmZmZmZmZmZERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVEREQzMzMzMzNVVVVVVVVmZmZ3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3dmZmZVVVVERERERERmZmZ3d3eIiIh3d3d3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZ3d3d3d3eIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVERERVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVERERERERERERVVVVVVVVERERERERERERERERVVVVVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZ3d3d3d3dmZmZmZmZmZmZmZmZ3d3d3d3dmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3dmZmZmZmZ3d3dmZmZVVVVmZmZmZmZ3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZEREREREQzMzNERERVVVVVVVUzMzNERERERERVVVVEREREREREREREREREREREREREREQzMzNEREREREREREREREREREREREREREREREREREREREQzMzNEREREREREREREREQzMzNERERVVVVERERVVVVEREREREREREREREREREQzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNEREQzMzMzMzNERERVVVVERERVVVVmZmZmZmZVVVVEREQzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzNEREREREQzMzMiIiIiIiIzMzMzMzNEREREREREREREREREREREREREREREREREREREREREREREREREREQzMzMzMzNEREQzMzNEREREREREREREREQzMzNERERVVVVVVVVEREREREREREREREREREQzMzNERERVVVVERERERERERERVVVVVVVVmZmZVVVVEREREREREREQzMzMzMzMzMzNEREREREQzMzN3d3eZmZlmZmZVVVVmZmZmZmZ3d3d3d3d3d3dVVVVEREREREREREREREREREREREQzMzMzMzNEREREREREREQzMzNERERmZmZEREREREQzMzNERERERERmZmaZmZmqqqqZmZmIiIiIiIiIiIhmZmZVVVVmZmZmZmZVVVVERERERERVVVVmZmZVVVVVVVVERERERERERERERERmZmZmZmZmZmZVVVVmZmZmZmZVVVVVVVVERERERERVVVVEREREREQzMzNEREREREQzMzMiIiIzMzMzMzMzMzMzMzNEREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERVVVVVVVVVVVVVVVVEREQzMzMzMzNERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERERERVVVV3d3eIiIh3d3eIiIiqqqqZmZmIiIiIiIh3d3eIiIiIiIh3d3dmZmZVVVUzMzNVVVWIiIiIiIhmZmZVVVVVVVVVVVVERERVVVVEREQzMzNEREREREQzMzNERERVVVVmZmaIiIiIiIh3d3dVVVVERERVVVV3d3d3d3dVVVUzMzMzMzMzMzMzMzNERERERERERERERERERERERERERERERERmZmZ3d3dmZmZVVVVmZmZVVVVERERERERERERERERERERERERVVVVVVVVVVVVVVVVmZmZ3d3dmZmZVVVVVVVVERERERERVVVVVVVVERERmZmZ3d3dmZmZVVVVmZmZ3d3dVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVV3d3d3d3d3d3dmZmZVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZVVVVmZmaIiIiZmZmIiIhVVVVVVVVmZmZmZmZmZmZmZmZ3d3eIiIh3d3eIiIiZmZl3d3dmZmZVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3dVVVVVVVVVVVVVVVVmZmZEREQzMzNERER3d3eIiIiIiIhmZmZmZmZVVVVERERERERVVVVmZmZmZmZmZmZmZmZmZmZ3d3eIiIiIiIi7u7uqqqqqqqrd3d3d3d3u7u7d3d27u7uIiIiIiIiIiIiIiIiIiIiIiIiZmZmIiIiIiIiZmZmZmZmZmZmIiIiZmZnMzMzMzMy7u7u7u7u7u7uqqqrMzMzMzMzMzMzMzMzd3d3////////////////u7u7///////////////////////////8A////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////7u7u////////////7u7u7u7u3d3dzMzMzMzMu7u7mZmZmZmZiIiIqqqqqqqqqqqqqqqqmZmZmZmZqqqqqqqqmZmZqqqqqqqqqqqqu7u7zMzMzMzMzMzMzMzMu7u7u7u7u7u7zMzMzMzMzMzMu7u7zMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7u7u7u7u7qqqqqqqqu7u7qqqqqqqqqqqqqqqqqqqqqqqqmZmZmZmZiIiImZmZiIiIiIiIiIiIiIiIiIiIiIiImZmZiIiIiIiIiIiImZmZiIiImZmZiIiIiIiId3d3iIiIiIiId3d3iIiIiIiIiIiIiIiId3d3iIiId3d3iIiId3d3iIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3iIiId3d3iIiId3d3d3d3iIiId3d3iIiIiIiIiIiId3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3iIiId3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmd3d3d3d3ZmZmd3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3ZmZmVVVVZmZmd3d3VVVVVVVVVVVVREREVVVVVVVVZmZmZmZmZmZmVVVVZmZmVVVVZmZmZmZmd3d3d3d3iIiIiIiIiIiImZmZmZmZd3d3iIiImZmZmZmZmZmZmZmZiIiIiIiId3d3iIiId3d3d3d3iIiImZmZiIiIiIiImZmZiIiId3d3iIiId3d3ZmZmVVVVVVVVu7u77u7uzMzMzMzMzMzM3d3dzMzMqqqqqqqqu7u7zMzMu7u7mZmZiIiImZmZqqqqu7u7qqqqqqqqqqqqmZmZqqqqqqqqqqqqiIiIZmZmZmZmd3d3iIiImZmZmZmZiIiIZmZmZmZmd3d3mZmZiIiIiIiIiIiIiIiId3d3iIiIiIiIiIiId3d3ZmZmVVVVREREmZmZqqqqmZmZmZmZmZmZiIiIiIiIiIiImZmZd3d3iIiImZmZmZmZmZmZiIiId3d3d3d3ZmZmiIiIiIiImZmZmZmZiIiIiIiId3d3ZmZmZmZmZmZmiIiId3d3iIiId3d3ZmZmd3d3d3d3VVVVVVVVd3d3ZmZmd3d3iIiImZmZiIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmVVVVVVVVVVVVZmZmd3d3d3d3iIiIiIiId3d3d3d3d3d3ZmZmiIiId3d3d3d3ZmZmVVVVVVVVREREREREVVVVVVVVd3d3iIiId3d3ZmZmZmZmd3d3ZmZmZmZmZmZmVVVVZmZmVVVVVVVVREREVVVVREREREREVVVVZmZmZmZmd3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmVVVVd3d3d3d3d3d3d3d3ZmZmREREVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVREREVVVVd3d3ZmZmd3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3iIiIZmZmVVVVVVVVZmZmZmZmd3d3REREVVVVVVVVVVVVVVVVZmZmZmZmd3d3iIiIiIiId3d3d3d3ZmZmREREREREREREREREVVVVZmZmZmZmVVVVVVVVZmZmVVVVVVVVREREVVVVVVVVZmZmZmZmZmZmVVVVZmZmREREREREMzMzVVVVZmZmd3d3ZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVZmZmd3d3d3d3ZmZmZmZmVVVVVVVVZmZmZmZmd3d3d3d3d3d3ZmZmVVVVVVVVVVVVZmZmVVVVVVVVVVVVZmZmd3d3iIiIiIiIiIiIiIiId3d3d3d3d3d3iIiIiIiId3d3d3d3ZmZmZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREREREVVVVVVVVZmZmZmZmZmZmd3d3ZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmd3d3ZmZmd3d3d3d3d3d3d3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmZmZmd3d3d3d3ZmZmZmZmiIiId3d3d3d3d3d3ZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREREREMzMzMzMzREREREREMzMzMzMzMzMzREREMzMzREREREREREREREREREREREREREREREREVVVVVVVVREREREREREREREREREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREREREVVVVVVVVVVVVVVVVVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREREREREREVVVVREREVVVVREREREREREREREREREREMzMzREREMzMzREREREREREREREREREREMzMzREREREREREREVVVVREREREREREREMzMzREREREREREREVVVVREREREREREREREREVVVVVVVVREREMzMzMzMzREREREREREREMzMzREREREREREREd3d3mZmZZmZmVVVVZmZmZmZmZmZmd3d3d3d3d3d3ZmZmVVVVREREREREMzMzREREREREMzMzREREMzMzREREMzMzMzMzVVVVREREMzMzMzMzREREVVVVVVVViIiImZmZmZmZiIiIiIiIiIiIZmZmREREZmZmVVVVZmZmREREREREREREVVVVZmZmVVVVVVVVVVVVREREZmZmZmZmd3d3ZmZmVVVVVVVVVVVVZmZmZmZmZmZmVVVVREREREREMzMzMzMzREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzREREMzMzMzMzREREMzMzMzMzMzMzREREMzMzMzMzREREVVVVVVVVVVVVVVVVREREMzMzREREMzMzREREREREREREVVVVVVVVVVVVREREREREREREREREREREREREREREVVVVd3d3iIiId3d3d3d3mZmZmZmZiIiIiIiIiIiIiIiId3d3ZmZmZmZmZmZmREREVVVViIiIiIiIZmZmZmZmVVVVVVVVREREREREREREMzMzREREREREREREREREVVVVREREVVVVZmZmVVVVVVVVREREVVVVd3d3iIiIZmZmREREMzMzMzMzMzMzMzMzMzMzREREMzMzVVVVREREREREVVVVVVVVVVVVZmZmVVVVVVVVVVVVZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVZmZmVVVVZmZmVVVVZmZmd3d3ZmZmVVVVVVVVVVVVREREVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3VVVVVVVVZmZmZmZmZmZmVVVVREREVVVVd3d3ZmZmVVVVVVVVZmZmVVVVVVVVd3d3iIiIiIiId3d3ZmZmZmZmd3d3d3d3ZmZmREREd3d3iIiId3d3iIiIiIiId3d3VVVVVVVVZmZmd3d3iIiId3d3d3d3iIiId3d3ZmZmZmZmVVVVVVVVVVVVMzMzMzMzVVVVmZmZmZmZmZmZZmZmVVVVVVVVZmZmVVVVZmZmZmZmVVVVVVVVZmZmZmZmd3d3d3d3d3d3iIiImZmZmZmZqqqqzMzMu7u7u7u7iIiIZmZmZmZmd3d3d3d3d3d3iIiImZmZiIiIiIiIqqqqmZmZiIiIiIiIiIiIqqqqqqqqqqqqqqqqqqqqqqqqu7u7u7u7zMzMzMzM7u7u////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7szMzLu7u6qqqpmZmZmZmaqqqszMzMzMzMzMzMzMzMzMzMzMzN3d3d3d3czMzN3d3d3d3e7u7t3d3e7u7u7u7u7u7u7u7t3d3e7u7u7u7u7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u6qqqru7u6qqqqqqqqqqqqqqqpmZmZmZmaqqqpmZmaqqqqqqqpmZmZmZmZmZmZmZmYiIiIiIiJmZmYiIiJmZmZmZmYiIiIiIiJmZmYiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d2ZmZoiIiHd3d3d3d2ZmZmZmZnd3d2ZmZmZmZnd3d3d3d3d3d2ZmZnd3d2ZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZnd3d2ZmZnd3d2ZmZnd3d4iIiHd3d3d3d4iIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d2ZmZmZmZmZmZnd3d4iIiIiIiHd3d3d3d4iIiHd3d2ZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVURERGZmZlVVVVVVVVVVVVVVVWZmZnd3d4iIiGZmZmZmZnd3d3d3d3d3d4iIiIiIiIiIiJmZmZmZmZmZmZmZmYiIiIiIiIiIiGZmZmZmZmZmZmZmZnd3d4iIiJmZmYiIiIiIiIiIiIiIiHd3d3d3d3d3d0RERERERGZmZru7u8zMzMzMzLu7u7u7u8zMzMzMzLu7u8zMzMzMzMzMzKqqqoiIiIiIiJmZmZmZmaqqqqqqqpmZmaqqqqqqqpmZmZmZmZmZmXd3d3d3d2ZmZnd3d5mZmZmZmYiIiIiIiHd3d2ZmZnd3d4iIiIiIiIiIiJmZmYiIiIiIiIiIiHd3d3d3d2ZmZmZmZlVVVVVVVYiIiJmZmYiIiJmZmZmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiJmZmZmZmXd3d2ZmZmZmZmZmZoiIiHd3d3d3d4iIiIiIiHd3d2ZmZmZmZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVVVVVWZmZlVVVWZmZnd3d3d3d2ZmZmZmZmZmZnd3d2ZmZmZmZmZmZnd3d3d3d2ZmZmZmZmZmZlVVVURERFVVVWZmZnd3d4iIiHd3d3d3d3d3d3d3d2ZmZnd3d4iIiHd3d3d3d1VVVVVVVURERERERERERERERFVVVWZmZnd3d2ZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZnd3d2ZmZlVVVVVVVVVVVURERERERFVVVVVVVWZmZmZmZmZmZmZmZnd3d3d3d4iIiHd3d3d3d3d3d3d3d2ZmZnd3d2ZmZlVVVVVVVWZmZnd3d2ZmZmZmZmZmZlVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZkRERFVVVVVVVXd3d3d3d3d3d3d3d2ZmZnd3d2ZmZnd3d4iIiHd3d3d3d3d3d4iIiHd3d2ZmZkRERFVVVWZmZmZmZnd3d1VVVVVVVURERFVVVWZmZlVVVWZmZnd3d3d3d4iIiIiIiIiIiHd3d2ZmZlVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVURERFVVVXd3d3d3d2ZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d5mZmXd3d3d3d2ZmZnd3d2ZmZmZmZlVVVVVVVVVVVWZmZnd3d4iIiIiIiJmZmZmZmZmZmZmZmYiIiHd3d2ZmZnd3d4iIiHd3d3d3d2ZmZmZmZmZmZmZmZnd3d3d3d2ZmZnd3d2ZmZlVVVVVVVWZmZmZmZlVVVXd3d3d3d3d3d2ZmZmZmZmZmZmZmZnd3d2ZmZmZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZnd3d2ZmZlVVVVVVVWZmZlVVVVVVVVVVVURERFVVVWZmZlVVVVVVVVVVVVVVVVVVVWZmZnd3d2ZmZmZmZlVVVWZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZlVVVVVVVWZmZmZmZmZmZmZmZmZmZnd3d3d3d4iIiHd3d2ZmZnd3d3d3d2ZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZmZmZmZmZmZmZnd3d3d3d2ZmZnd3d4iIiGZmZlVVVURERERERDMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM0RERDMzMzMzM0RERERERDMzM0RERFVVVURERFVVVURERFVVVVVVVVVVVVVVVURERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERERERFVVVVVVVURERFVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERERERERERDMzM0RERDMzM0RERDMzM0RERERERERERFVVVURERERERERERERERDMzM0RERDMzM0RERERERFVVVURERDMzM0RERDMzM0RERDMzM0RERERERERERDMzM0RERERERFVVVVVVVURERERERFVVVURERERERERERERERERERDMzMzMzM0RERFVVVVVVVVVVVVVVVVVVVURERFVVVWZmZmZmZlVVVWZmZmZmZnd3d3d3d2ZmZnd3d2ZmZlVVVURERERERERERERERERERERERERERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVWZmZoiIiJmZmZmZmZmZmXd3d2ZmZmZmZlVVVWZmZmZmZlVVVURERFVVVURERFVVVURERFVVVVVVVVVVVURERGZmZnd3d3d3d3d3d2ZmZmZmZnd3d2ZmZmZmZnd3d1VVVVVVVTMzMzMzMzMzMzMzM0RERERERERERCIiIjMzMzMzMzMzM0RERDMzMzMzM0RERERERDMzMzMzMzMzMyIiIjMzMzMzMzMzM1VVVVVVVVVVVVVVVURERERERDMzMzMzM0RERERERERERERERFVVVVVVVVVVVVVVVVVVVURERERERERERERERERERFVVVXd3d4iIiGZmZmZmZnd3d4iIiIiIiHd3d3d3d4iIiJmZmYiIiHd3d3d3d0RERERERIiIiIiIiGZmZmZmZlVVVVVVVURERERERERERERERERERERERERERERERERERERERERERFVVVVVVVVVVVURERFVVVVVVVWZmZnd3d1VVVURERDMzMzMzMzMzM0RERDMzM0RERERERERERERERERERFVVVURERFVVVVVVVURERGZmZnd3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVURERERERFVVVWZmZmZmZnd3d2ZmZlVVVVVVVWZmZlVVVVVVVURERGZmZnd3d1VVVVVVVVVVVVVVVWZmZnd3d3d3d4iIiIiIiIiIiJmZmZmZmZmZmYiIiGZmZlVVVWZmZnd3d3d3d2ZmZmZmZmZmZnd3d2ZmZnd3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiGZmZmZmZmZmZlVVVTMzMzMzM1VVVaqqqru7u5mZmXd3d1VVVWZmZmZmZnd3d2ZmZmZmZmZmZlVVVVVVVXd3d2ZmZmZmZmZmZmZmZnd3d3d3d3d3d4iIiJmZmYiIiGZmZnd3d2ZmZmZmZmZmZnd3d3d3d4iIiJmZmYiIiJmZmZmZmZmZmaqqqpmZmaqqqqqqqqqqqqqqqru7u6qqqru7u7u7u7u7u8zMzP///////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////u7u7////////////////////////////u7u7u7u7u7u7////u7u7////////u7u7u7u7u7u7u7u7u7u7d3d3d3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7d3d3d3d3d3d3d3d3MzMzMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3MzMzd3d3MzMzMzMzMzMzMzMy7u7vMzMy7u7vMzMy7u7u7u7u7u7u7u7uqqqq7u7uqqqqqqqq7u7uqqqqqqqqZmZmqqqqZmZmIiIiZmZmIiIiIiIiIiIiIiIh3d3d3d3d3d3dmZmZ3d3d3d3dmZmZVVVVmZmZmZmZVVVVVVVV3d3dmZmZmZmZ3d3dmZmZ3d3dmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3eIiIiIiIiIiIiIiIiZmZmIiIiZmZmZmZmZmZmZmZmZmZmIiIiZmZmZmZmIiIiZmZmIiIiZmZmIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZ3d3d3d3eZmZmqqqqZmZlmZmZmZmZ3d3d3d3eZmZmZmZmIiIiZmZmIiIiIiIh3d3eIiIh3d3d3d3dVVVVVVVVmZmZVVVV3d3eZmZmZmZmIiIh3d3d3d3eIiIiIiIiIiIhmZmZVVVVVVVVmZma7u7vd3d27u7uqqqqqqqqqqqrMzMzMzMzMzMzd3d3d3d2qqqqZmZmIiIiZmZmqqqqZmZmqqqqqqqqqqqqqqqqZmZmZmZmZmZmIiIh3d3dmZmZ3d3eIiIiIiIh3d3d3d3dmZmZmZmZ3d3eIiIiIiIiZmZmZmZmIiIiIiIiIiIh3d3d3d3d3d3dmZmZERERERESIiIiIiIh3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiZmZmZmZmIiIiIiIh3d3d3d3dmZmZVVVV3d3dVVVV3d3eZmZmIiIh3d3dmZmZ3d3d3d3eIiIh3d3dmZmZmZmZmZmZmZmZmZmZmZmZVVVVERERVVVVERERVVVV3d3dmZmZmZmZmZmZVVVVmZmZmZmZVVVV3d3d3d3dmZmZ3d3dmZmZVVVVERERVVVVVVVVVVVVmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3d3d3dVVVVERERVVVVERERVVVVERERERERVVVVmZmaIiIh3d3dmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVERERERERVVVVmZmZmZmZ3d3dmZmZmZmZ3d3d3d3eIiIh3d3eIiIh3d3dmZmZmZmZmZmZVVVVERERVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVV3d3dVVVVVVVVVVVVVVVVmZmZ3d3d3d3d3d3dmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3eIiIh3d3dmZmZVVVVVVVVmZmZ3d3eIiIhmZmZVVVVERERVVVVVVVVmZmZmZmZ3d3d3d3d3d3eIiIiIiIiIiIh3d3d3d3d3d3eIiIh3d3d3d3d3d3dVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZ3d3d3d3d3d3dmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmaIiIiqqqqqqqqZmZmIiIiZmZmZmZmIiIh3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIiqqqqZmZl3d3d3d3dmZmZ3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZ3d3eIiIhmZmZmZmZmZmZVVVVmZmZmZmZ3d3dmZmZVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZVVVVVVVVVVVVVVVVERERVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3dVVVVmZmZ3d3dmZmaIiIiIiIh3d3dmZmZ3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3dmZmZmZmZVVVVVVVVmZmZmZmZVVVVmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIhmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVEREREREQzMzNEREQzMzMzMzMzMzMzMzNERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzNERERERERERERERERVVVVERERERERERERVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzNERERERERVVVVEREREREREREREREREREREREREREREREREREQzMzNERERVVVVERERVVVVERERERERERERERERERERERERERERVVVVEREREREREREREREREREQzMzMzMzMzMzNERERERERERERERERERERmZmZVVVVERERVVVVEREREREQzMzMzMzMzMzNEREREREQzMzMzMzNERERVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3dVVVVEREREREREREREREREREQzMzNEREREREQzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNVVVVVVVV3d3eZmZmZmZmIiIh3d3dmZmZVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVERERERERERERVVVVVVVVERERmZmaIiIh3d3dmZmZVVVVVVVVmZmZmZmZmZmZ3d3dmZmZVVVVEREREREQzMzNERERERERVVVUzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVEREQzMzMiIiJEREREREQzMzNEREREREREREREREREREREREREREREREREREQzMzNERERERERERERERERVVVVVVVVVVVVVVVVEREQzMzMzMzNERERERERVVVVmZmZ3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmaIiIiqqqqZmZmqqqpmZmZERER3d3eIiIhmZmZVVVVVVVVVVVVVVVVEREREREREREQzMzNERERERERERERERERERERERERERERERERVVVVVVVVERERVVVVVVVVmZmZ3d3dVVVUzMzMzMzMzMzMzMzNEREQzMzNERERERERERERVVVVERERVVVVERERERERVVVVVVVVmZmZVVVVERERVVVVVVVVERERVVVVERERVVVVERERVVVVVVVVVVVVERERVVVVmZmZ3d3dmZmZmZmZVVVVVVVVVVVVmZmZVVVVVVVVVVVVERERERERVVVVERERERERVVVVmZmZmZmZERERVVVVmZmZVVVVVVVVVVVVmZmZ3d3d3d3dmZmZmZmZmZmZ3d3eZmZmIiIiIiIiqqqq7u7u7u7uqqqqZmZmIiIh3d3dVVVVVVVVmZmZ3d3dmZmZmZmZmZmZmZmaIiIhmZmZmZmZ3d3d3d3eZmZmqqqqZmZmIiIhmZmZmZmZ3d3dVVVVEREQzMzNERESZmZnMzMyqqqp3d3dVVVVmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZ3d3d3d3dmZmZmZmZmZmZ3d3eIiIh3d3d3d3eIiIh3d3eIiIh3d3eIiIiIiIiZmZmIiIiqqqqIiIiZmZmqqqqqqqqqqqq7u7uqqqqqqqq7u7u7u7u7u7u7u7u7u7u7u7vd3d3u7u7///////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzM3d3dzMzM3d3d3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7zMzMu7u7qqqqqqqqqqqqmZmZmZmZmZmZiIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZiIiImZmZiIiIiIiIiIiImZmZmZmZmZmZqqqqqqqqmZmZmZmZqqqqqqqqmZmZmZmZmZmZmZmZqqqqqqqqqqqqmZmZqqqqmZmZiIiIiIiIiIiImZmZiIiIiIiIiIiImZmZiIiImZmZiIiIiIiIiIiId3d3d3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVVVVVREREREREVVVVREREVVVVREREVVVVREREVVVVREREVVVVVVVVd3d3iIiId3d3d3d3d3d3iIiId3d3iIiIqqqqu7u7zMzMmZmZZmZmZmZmd3d3d3d3d3d3iIiId3d3ZmZmd3d3iIiIiIiId3d3ZmZmVVVVd3d3d3d3ZmZmd3d3iIiIiIiId3d3ZmZmZmZmd3d3iIiImZmZd3d3ZmZmVVVVd3d3u7u7zMzMu7u7u7u7u7u7u7u7u7u7u7u7zMzM3d3dzMzMqqqqiIiImZmZqqqqmZmZqqqqu7u7qqqqqqqqqqqqqqqqmZmZiIiId3d3d3d3ZmZmZmZmd3d3d3d3iIiId3d3ZmZmVVVVZmZmd3d3iIiImZmZmZmZmZmZiIiId3d3iIiId3d3ZmZmZmZmVVVVVVVVZmZmZmZmd3d3iIiId3d3d3d3iIiImZmZiIiIiIiImZmZmZmZd3d3d3d3iIiId3d3VVVVZmZmd3d3VVVVd3d3qqqqmZmZd3d3d3d3d3d3d3d3d3d3iIiIiIiId3d3VVVVVVVVVVVVZmZmVVVVVVVVREREREREVVVVZmZmZmZmZmZmd3d3ZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREVVVVd3d3d3d3d3d3d3d3ZmZmZmZmZmZmd3d3d3d3d3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVd3d3iIiIZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVREREVVVVVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmd3d3ZmZmVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3VVVVVVVVVVVVZmZmZmZmd3d3d3d3ZmZmVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3iIiIZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3VVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3iIiIiIiIiIiIZmZmd3d3mZmZd3d3ZmZmd3d3ZmZmVVVVREREVVVVREREVVVVZmZmZmZmZmZmZmZmVVVVZmZmVVVVZmZmd3d3d3d3iIiId3d3d3d3ZmZmVVVVZmZmVVVVVVVVVVVVVVVVZmZmREREVVVVZmZmVVVVVVVVZmZmd3d3iIiImZmZmZmZiIiId3d3d3d3d3d3d3d3d3d3ZmZmZmZmVVVVVVVVZmZmVVVVVVVVVVVVVVVVZmZmZmZmd3d3iIiId3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmd3d3iIiId3d3iIiId3d3d3d3d3d3ZmZmVVVVZmZmd3d3ZmZmVVVVVVVVVVVVVVVVREREREREREREVVVVREREREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVZmZmVVVVREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3ZmZmd3d3iIiId3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3ZmZmZmZmZmZmVVVVZmZmd3d3ZmZmZmZmd3d3d3d3d3d3d3d3ZmZmVVVVVVVVZmZmZmZmVVVVREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3iIiId3d3iIiIiIiId3d3d3d3d3d3ZmZmZmZmZmZmd3d3d3d3ZmZmd3d3ZmZmVVVVVVVVVVVVVVVVVVVVREREREREREREREREVVVVREREVVVVVVVVVVVVREREVVVVREREREREREREREREMzMzMzMzMzMzMzMzREREMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREMzMzREREREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzREREREREMzMzMzMzMzMzMzMzMzMzREREREREVVVVREREREREREREREREREREREREREREREREREREMzMzMzMzREREVVVVVVVVREREREREMzMzMzMzREREREREVVVVVVVVREREREREMzMzMzMzMzMzMzMzREREMzMzREREREREREREREREZmZmVVVVREREREREREREREREREREMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzREREREREMzMzREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3iIiId3d3d3d3ZmZmVVVVVVVVREREREREREREREREREREREREREREIiIiMzMzIiIiMzMzIiIiMzMzMzMzREREVVVVZmZmiIiImZmZiIiIZmZmZmZmZmZmVVVVVVVVVVVVd3d3ZmZmZmZmVVVVREREREREREREREREVVVVREREVVVVd3d3VVVVREREVVVVVVVVVVVVZmZmZmZmZmZmVVVVREREREREREREVVVVVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzZmZmVVVVMzMzMzMzREREREREVVVVREREREREREREREREREREREREREREREREREREREREREREREREVVVVVVVVREREZmZmZmZmVVVVREREREREMzMzREREREREVVVVZmZmZmZmd3d3d3d3d3d3d3d3ZmZmd3d3VVVVZmZmiIiImZmZqqqqu7u7ZmZmMzMzZmZmd3d3VVVVVVVVREREREREREREREREVVVVREREMzMzREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVREREVVVVZmZmd3d3d3d3ZmZmREREMzMzREREMzMzREREMzMzREREREREVVVVREREREREREREREREREREVVVVREREREREREREREREREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVREREREREVVVVREREREREREREREREVVVVREREVVVVVVVVVVVVVVVVREREREREVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3ZmZmiIiIiIiIiIiIiIiId3d3mZmZqqqqmZmZd3d3iIiIiIiIVVVVVVVVZmZmd3d3ZmZmVVVVVVVVVVVVZmZmZmZmd3d3d3d3iIiImZmZqqqqiIiId3d3ZmZmd3d3d3d3VVVVVVVVMzMzREREiIiIu7u7u7u7iIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiId3d3iIiId3d3d3d3d3d3iIiIqqqqu7u7qqqqqqqqqqqqqqqqmZmZqqqqqqqqu7u73d3du7u7qqqqu7u7u7u7zMzMzMzMu7u7zMzM3d3d////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7t3d3d3d3e7u7t3d3d3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3e7u7u7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3czMzMzMzMzMzMzMzLu7u7u7u6qqqqqqqqqqqqqqqpmZmZmZmZmZmYiIiJmZmZmZmZmZmYiIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiIiIiIiIiIiIiJmZmZmZmZmZmZmZmYiIiIiIiIiIiIiIiIiIiJmZmYiIiKqqqpmZmaqqqpmZmZmZmZmZmZmZmaqqqpmZmaqqqpmZmaqqqpmZmaqqqqqqqpmZmaqqqqqqqpmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiIiIiJmZmYiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERERERDMzM0RERFVVVURERFVVVVVVVURERFVVVWZmZlVVVWZmZmZmZnd3d4iIiIiIiHd3d2ZmZnd3d2ZmZmZmZoiIiLu7u93d3d3d3bu7u3d3d2ZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZoiIiIiIiHd3d3d3d3d3d4iIiIiIiHd3d4iIiIiIiGZmZnd3d2ZmZlVVVWZmZnd3d4iIiHd3d3d3d2ZmZoiIiLu7u8zMzMzMzMzMzKqqqru7u8zMzLu7u8zMzMzMzMzMzLu7u6qqqpmZmaqqqpmZmaqqqqqqqqqqqqqqqqqqqpmZmZmZmYiIiHd3d3d3d2ZmZmZmZmZmZoiIiIiIiGZmZmZmZlVVVWZmZnd3d3d3d4iIiIiIiJmZmZmZmYiIiIiIiHd3d2ZmZmZmZlVVVURERFVVVXd3d3d3d4iIiIiIiHd3d3d3d4iIiJmZmYiIiIiIiIiIiIiIiIiIiHd3d2ZmZlVVVWZmZmZmZlVVVWZmZpmZmZmZmYiIiHd3d3d3d3d3d2ZmZnd3d3d3d3d3d2ZmZlVVVWZmZlVVVVVVVURERERERERERFVVVWZmZmZmZmZmZnd3d2ZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZlVVVWZmZnd3d1VVVVVVVVVVVXd3d3d3d3d3d3d3d2ZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZlVVVVVVVWZmZmZmZlVVVVVVVWZmZmZmZnd3d2ZmZlVVVVVVVWZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZnd3d2ZmZnd3d2ZmZlVVVVVVVWZmZmZmZlVVVVVVVURERFVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZnd3d3d3d2ZmZmZmZlVVVWZmZlVVVWZmZnd3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d3d3d3d3d4iIiHd3d3d3d2ZmZmZmZlVVVVVVVWZmZlVVVWZmZmZmZmZmZnd3d3d3d4iIiIiIiHd3d3d3d4iIiHd3d2ZmZmZmZnd3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVWZmZnd3d3d3d2ZmZnd3d3d3d2ZmZlVVVVVVVVVVVVVVVWZmZmZmZnd3d1VVVVVVVVVVVWZmZmZmZnd3d3d3d4iIiHd3d3d3d4iIiHd3d2ZmZmZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVURERFVVVVVVVURERFVVVVVVVWZmZnd3d2ZmZmZmZlVVVWZmZmZmZlVVVVVVVWZmZmZmZlVVVWZmZmZmZmZmZnd3d3d3d2ZmZlVVVWZmZlVVVWZmZmZmZnd3d4iIiIiIiIiIiHd3d3d3d2ZmZmZmZnd3d2ZmZnd3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVURERFVVVVVVVURERFVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVURERFVVVVVVVVVVVWZmZmZmZnd3d3d3d3d3d2ZmZnd3d3d3d3d3d4iIiHd3d4iIiHd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZnd3d3d3d2ZmZmZmZmZmZnd3d2ZmZlVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d3d3d3d3d4iIiIiIiHd3d3d3d3d3d3d3d2ZmZmZmZlVVVWZmZnd3d2ZmZmZmZmZmZmZmZnd3d2ZmZlVVVWZmZlVVVVVVVWZmZlVVVWZmZlVVVVVVVURERERERDMzM0RERERERDMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERDMzM0RERDMzM0RERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzM0RERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERFVVVURERERERERERERERERERFVVVURERFVVVURERERERERERDMzM0RERERERDMzM0RERERERERERFVVVVVVVWZmZlVVVVVVVURERERERERERDMzMzMzMzMzMzMzM0RERDMzM0RERDMzMyIiIjMzM0RERDMzMzMzM0RERFVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d3d3d3d3d3d3d3d3d2ZmZlVVVURERERERERERFVVVURERFVVVURERDMzMzMzMzMzMyIiIjMzMyIiIiIiIjMzM1VVVWZmZoiIiJmZmZmZmYiIiHd3d3d3d2ZmZkRERFVVVXd3d3d3d2ZmZlVVVVVVVVVVVURERERERFVVVVVVVVVVVWZmZlVVVVVVVVVVVURERFVVVVVVVWZmZlVVVURERERERERERFVVVWZmZlVVVURERERERDMzM0RERDMzMzMzMzMzMzMzM0RERDMzMyIiIkRERFVVVURERERERDMzM0RERFVVVVVVVTMzMzMzM0RERERERERERERERDMzM0RERERERERERERERERERERERERERFVVVVVVVVVVVURERERERDMzM0RERERERFVVVVVVVVVVVXd3d2ZmZmZmZmZmZnd3d2ZmZlVVVVVVVYiIiJmZmaqqqru7u2ZmZjMzM2ZmZnd3d2ZmZlVVVURERERERFVVVURERFVVVURERERERDMzMzMzM0RERERERERERERERERERFVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVXd3d3d3d2ZmZlVVVURERERERERERDMzM0RERERERERERFVVVVVVVURERFVVVVVVVVVVVURERERERERERERERFVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVURERFVVVVVVVVVVVVVVVWZmZlVVVVVVVURERERERERERERERERERFVVVVVVVVVVVWZmZmZmZlVVVWZmZmZmZlVVVVVVVURERFVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d3d3d4iIiGZmZnd3d3d3d4iIiIiIiGZmZmZmZmZmZmZmZlVVVURERGZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZoiIiIiIiHd3d4iIiJmZmYiIiHd3d4iIiHd3d2ZmZmZmZmZmZkRERDMzM1VVVZmZmaqqqoiIiHd3d3d3d3d3d4iIiHd3d4iIiIiIiHd3d4iIiIiIiIiIiIiIiIiIiJmZmYiIiIiIiIiIiJmZmXd3d4iIiIiIiGZmZmZmZlVVVXd3d5mZmaqqqru7u6qqqru7u6qqqqqqqqqqqru7u8zMzMzMzLu7u7u7u6qqqru7u8zMzMzMzN3d3d3d3f///////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7d3d3u7u7u7u7u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzd3d3MzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7uqqqq7u7u7u7uqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqZmZmqqqqZmZmZmZmZmZmZmZmIiIiZmZmqqqqZmZmZmZmZmZmqqqqqqqqZmZmZmZmZmZmZmZmqqqqqqqqqqqqqqqqqqqqZmZmqqqqqqqqZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmIiIiIiIiIiIiZmZmIiIiIiIh3d3d3d3d3d3dmZmZVVVV3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVERERmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZ3d3eIiIh3d3d3d3eIiIhmZmZmZmZ3d3dVVVVmZmaZmZnMzMzd3d3d3d2qqqqIiIh3d3dVVVV3d3d3d3dmZmZ3d3eIiIh3d3dmZmaIiIh3d3eIiIiZmZmZmZmZmZl3d3d3d3d3d3dVVVVmZmZVVVVVVVVmZmZmZmZmZmZ3d3eIiIhmZmZ3d3e7u7vMzMzMzMy7u7uqqqqqqqqqqqq7u7vMzMzMzMzd3d2qqqqZmZmZmZmIiIiIiIiZmZmqqqqqqqqqqqqqqqqqqqqIiIiZmZl3d3dmZmZVVVVVVVV3d3d3d3eIiIiIiIh3d3dVVVVmZmZ3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIh3d3dmZmZmZmZVVVVERERVVVWIiIiIiIh3d3d3d3d3d3eIiIiIiIiIiIiIiIiZmZmIiIiIiIiIiIhmZmZVVVVmZmaIiIh3d3dmZmZ3d3eZmZmZmZmIiIiIiIh3d3dmZmZmZmZmZmZ3d3dVVVVmZmZmZmZVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3dmZmZVVVVVVVVmZmZ3d3dVVVVVVVVmZmZ3d3eIiIh3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmaIiIh3d3dmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZmZmZVVVVmZmZmZmZmZmZmZmZ3d3eIiIiIiIiIiIhmZmZmZmZ3d3d3d3dmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3eIiIhmZmZVVVVmZmZ3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZ3d3d3d3eIiIh3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZ3d3d3d3eIiIiIiIiIiIiZmZmZmZmZmZmZmZl3d3dmZmZ3d3d3d3dmZmZVVVVVVVVmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3eZmZmZmZmZmZmIiIiIiIh3d3d3d3d3d3d3d3dmZmZmZmZmZmZVVVVVVVVmZmZmZmZVVVVVVVVmZmZ3d3d3d3dmZmZ3d3d3d3dmZmZVVVVVVVVERERVVVVmZmZ3d3eZmZmqqqqIiIiIiIiIiIiIiIiZmZmZmZmZmZmIiIh3d3d3d3d3d3dVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVERERERERVVVVVVVVmZmZmZmZVVVVmZmZmZmZmZmZ3d3dmZmZmZmZVVVVmZmZ3d3dmZmZVVVVmZmaIiIh3d3d3d3dmZmZVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZVVVVERERVVVVERERERERVVVVVVVVVVVVmZmZVVVVmZmZVVVVmZmZ3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIhmZmZVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3dVVVVmZmZVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3dmZmZmZmZVVVVVVVVmZmZVVVVmZmZmZmZVVVVmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZmZmYA//8AAFVVVVVVVVVVVVVVVURERERERDMzM0RERFVVVURERDMzMyIiIiIiIjMzMyIiIiIiIjMzMzMzMzMzM0RERERERERERERERFVVVVVVVVVVVTMzMzMzMzMzMzMzMzMzM0RERERERERERERERDMzM0RERERERDMzMzMzMzMzMyIiIjMzM0RERERERERERERERERERERERERERERERERERDMzM0RERERERERERERERDMzM0RERERERERERDMzMzMzM0RERERERFVVVVVVVURERERERERERERERERERERERDMzM0RERERERFVVVURERERERGZmZmZmZkRERFVVVURERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMyIiIjMzMzMzM0RERERERERERFVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d1VVVVVVVURERFVVVVVVVVVVVVVVVURERDMzMzMzMyIiIjMzMyIiIjMzMzMzM0RERFVVVWZmZnd3d6qqqru7u5mZmXd3d3d3d2ZmZlVVVURERGZmZoiIiGZmZlVVVVVVVVVVVURERERERFVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVURERFVVVVVVVVVVVVVVVURERFVVVWZmZlVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERGZmZkRERDMzMzMzM1VVVURERDMzM0RERERERERERFVVVURERERERERERERERERERERERFVVVURERFVVVVVVVVVVVVVVVVVVVURERERERERERERERGZmZlVVVVVVVXd3d3d3d1VVVWZmZmZmZmZmZlVVVURERGZmZnd3d5mZmZmZmWZmZjMzM3d3d3d3d2ZmZlVVVVVVVURERERERFVVVVVVVURERERERERERERERERERERERERERDMzM1VVVVVVVWZmZmZmZnd3d2ZmZkRERERERFVVVXd3d4iIiIiIiGZmZlVVVTMzMzMzM0RERERERERERERERGZmZmZmZlVVVVVVVVVVVVVVVURERERERERERERERFVVVURERERERFVVVVVVVVVVVVVVVXd3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERFVVVURERFVVVVVVVWZmZnd3d2ZmZnd3d2ZmZnd3d2ZmZlVVVVVVVURERFVVVVVVVWZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZlVVVXd3d4iIiIiIiGZmZnd3d3d3d3d3d2ZmZkRERGZmZnd3d1VVVURERFVVVVVVVWZmZnd3d4iIiIiIiHd3d3d3d6qqqpmZmYiIiJmZmXd3d2ZmZoiIiIiIiGZmZkRERERERFVVVXd3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiJmZmYiIiJmZmYiIiIiIiJmZmYiIiIiIiJmZmZmZmYiIiKqqqpmZmWZmZlVVVVVVVVVVVXd3d5mZmaqqqszMzLu7u7u7u8zMzMzMzMzMzMzMzLu7u6qqqqqqqru7u8zMzMzMzMzMzO7u7v///////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////u7u7////////u7u7////u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7////u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3MzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7vMzMzMzMzd3d3MzMzMzMzd3d3MzMzd3d3MzMzd3d3d3d3MzMzd3d3MzMzMzMzMzMzMzMzMzMy7u7vMzMy7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7uqqqqqqqqqqqqZmZmZmZmqqqqZmZmqqqqZmZmZmZmIiIiZmZmZmZmIiIiIiIiZmZmZmZmqqqqqqqqqqqqqqqqZmZmZmZmZmZmZmZmZmZmIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIh3d3d3d3d3d3eIiIiIiIh3d3d3d3d3d3dmZmZ3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVVERERVVVVVVVVmZmZVVVVVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3dVVVVmZmZmZmZ3d3dmZmZmZmZmZmZVVVVVVVVmZmZVVVVmZmZVVVVmZmZ3d3dmZmZmZmZ3d3eZmZl3d3d3d3d3d3dmZmZ3d3d3d3d3d3eIiIiqqqqqqqq7u7uqqqqZmZmIiIhmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZ3d3d3d3eqqqq7u7uqqqqIiIhmZmZ3d3d3d3dmZmZVVVVVVVVVVVVERERVVVV3d3d3d3dVVVVVVVWqqqrMzMzMzMyqqqqZmZmqqqqIiIiqqqq7u7vMzMzMzMyqqqqZmZmIiIiZmZmZmZmIiIiZmZmqqqqqqqqqqqqZmZmZmZmIiIh3d3dVVVVERERERERmZmZ3d3eIiIiIiIh3d3dmZmZmZmZ3d3d3d3d3d3d3d3eIiIiIiIiIiIh3d3eIiIhmZmZVVVVERERERER3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiZmZmIiIiIiIh3d3d3d3dmZmZmZmaZmZmIiIh3d3dmZmZmZmaIiIiZmZmZmZmIiIh3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3dmZmZVVVVVVVVmZmZmZmZmZmZ3d3dVVVVmZmZVVVVmZmZmZmZ3d3dmZmZmZmZ3d3d3d3eIiIhmZmZVVVVmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZ3d3d3d3dmZmZmZmZ3d3dmZmZVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmaIiIiZmZmZmZmIiIh3d3d3d3d3d3dmZmZmZmZ3d3dmZmZmZmZVVVVmZmZVVVVmZmZ3d3d3d3eZmZmIiIiIiIh3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVmZmZmZmZmZmaIiIiIiIh3d3d3d3d3d3dmZmZVVVVmZmZmZmZmZmZVVVVmZmZVVVVmZmZmZmZmZmZ3d3eIiIiZmZmZmZmIiIiIiIh3d3dmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3eIiIiZmZmqqqqZmZmIiIiIiIh3d3d3d3dmZmZ3d3d3d3d3d3dmZmZVVVVVVVVmZmZmZmZVVVVmZmZ3d3d3d3dmZmZ3d3d3d3d3d3dmZmZmZmZVVVVERERVVVVVVVWIiIiqqqq7u7uZmZmZmZmZmZmZmZmqqqq7u7uZmZmIiIh3d3d3d3dmZmZVVVVmZmZVVVVmZmZVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVmZmZmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3dVVVVERERVVVVVVVVVVVVmZmZVVVVmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZVVVVERERVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVV3d3dmZmZmZmZmZmZVVVVmZmZVVVVmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZ3d3dmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3dmZmZ3d3eIiIhmZmZmZmaIiIhmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVERERVVVVVVVVVVVVmZmZVVVVmZmZVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZ3d3dmZmZ3d3d3d3dmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZVVVV3d3d3d3dmZmZVVVUzMzMzMzMiIiIzMzMiIiIzMzMiIiJEREREREREREREREREREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERVVVVEREREREREREQzMzMzMzNEREQzMzNERERERERERERERERVVVVERERERERERERERERERERVVVVERERERERERERVVVVEREREREREREREREREREQzMzNEREQzMzNERERVVVVmZmZVVVVVVVVERERVVVVEREQzMzMzMzMzMzMzMzMzMzNEREQzMzNEREREREREREQzMzMzMzMzMzNVVVVmZmZVVVVmZmZVVVVmZmZmZmZmZmZ3d3dmZmZmZmZ3d3d3d3d3d3dmZmZmZmZmZmZVVVVEREREREREREQzMzMzMzMzMzMiIiIiIiIzMzMzMzNERERERERVVVVVVVV3d3eqqqq7u7uqqqqIiIh3d3dmZmZVVVVERERVVVVVVVVmZmZVVVVmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVERERmZmZVVVVmZmZVVVVVVVVVVVVERERVVVVmZmZEREQzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMiIiIzMzNERERERERERERERERVVVVEREQzMzMzMzMzMzNVVVUzMzNEREREREREREREREREREREREREREQzMzNERERERERERERVVVVERERVVVVmZmZVVVVERERERERERERERERVVVVmZmZmZmZVVVV3d3dmZmZmZmZmZmZVVVVERERERERERERERERmZmZ3d3eIiIh3d3dERERmZmZ3d3dmZmZVVVVVVVVERERERERERERVVVVEREREREQzMzMzMzNERERERERVVVVERERERERVVVVVVVVmZmZ3d3dmZmZVVVVVVVVERERERER3d3e7u7uIiIhVVVVVVVVVVVVERERERERERERERERmZmZ3d3dmZmZmZmZVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVERERERERVVVVERERERERERERERERERERERERVVVVVVVVVVVVVVVVmZmZ3d3dmZmZ3d3d3d3dmZmZVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERmZmZ3d3eIiIiZmZmqqqqZmZmIiIh3d3dVVVVVVVVmZmZ3d3dmZmZmZmZmZmZ3d3eIiIiZmZm7u7uqqqqIiIiZmZm7u7u7u7uqqqqqqqp3d3eIiIiZmZmIiIh3d3dmZmZVVVVVVVV3d3d3d3dmZmZ3d3dmZmZmZmZmZmaIiIiZmZmZmZmIiIiIiIiIiIiZmZmIiIiIiIiIiIiZmZmqqqqqqqqIiIh3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3eIiIiqqqqqqqqqqqq7u7u7u7u7u7u7u7uZmZmZmZm7u7u7u7u7u7vMzMzd3d3///////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////7u7u////7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d7u7u7u7u3d3d3d3d7u7u3d3d3d3d3d3dzMzMzMzMzMzMu7u7u7u7qqqqu7u7qqqqu7u7u7u7zMzMzMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7u7u7qqqqu7u7qqqqqqqqmZmZmZmZmZmZmZmZiIiImZmZqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqmZmZmZmZmZmZmZmZmZmZmZmZd3d3d3d3d3d3iIiId3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmVVVVVVVVVVVVREREREREREREREREREREVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmd3d3ZmZmZmZmd3d3iIiIiIiId3d3ZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmd3d3ZmZmZmZmZmZmd3d3iIiIZmZmZmZmZmZmZmZmd3d3d3d3iIiImZmZmZmZmZmZqqqqmZmZd3d3d3d3d3d3d3d3iIiIiIiImZmZd3d3ZmZmd3d3iIiIiIiIiIiIqqqqqqqqmZmZd3d3ZmZmiIiIiIiIiIiId3d3ZmZmVVVVVVVViIiIiIiIiIiId3d3VVVVqqqq3d3dzMzMu7u7u7u7u7u7mZmZmZmZu7u7zMzMqqqqmZmZmZmZmZmZmZmZmZmZiIiImZmZmZmZmZmZqqqqmZmZmZmZmZmZd3d3ZmZmVVVVVVVVVVVViIiImZmZiIiId3d3d3d3ZmZmVVVVd3d3d3d3d3d3mZmZiIiIiIiId3d3d3d3ZmZmZmZmREREVVVVd3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiId3d3iIiIZmZmd3d3iIiIiIiIiIiId3d3ZmZmd3d3iIiImZmZd3d3ZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3iIiIiIiId3d3d3d3ZmZmVVVVVVVVd3d3d3d3d3d3ZmZmVVVVVVVVZmZmd3d3d3d3d3d3d3d3iIiImZmZiIiId3d3d3d3ZmZmZmZmZmZmd3d3d3d3VVVVVVVVZmZmZmZmd3d3ZmZmZmZmZmZmd3d3iIiIiIiId3d3d3d3ZmZmZmZmVVVVZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmiIiImZmZqqqqmZmZiIiId3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmiIiIiIiId3d3d3d3iIiIZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREVVVVREREVVVVZmZmVVVVZmZmd3d3iIiIiIiId3d3d3d3ZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmiIiIiIiIiIiIiIiIiIiId3d3ZmZmZmZmVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3iIiImZmZmZmZd3d3d3d3ZmZmZmZmZmZmVVVVd3d3d3d3d3d3ZmZmVVVVZmZmZmZmZmZmVVVVZmZmd3d3d3d3d3d3ZmZmd3d3ZmZmZmZmZmZmVVVVVVVVREREVVVVZmZmiIiId3d3ZmZmZmZmZmZmd3d3iIiIiIiIiIiId3d3d3d3ZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVREREREREVVVVd3d3ZmZmVVVVVVVVVVVVZmZmVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmd3d3ZmZmZmZmd3d3ZmZmd3d3d3d3d3d3ZmZmZmZmZmZmVVVVVVVVZmZmVVVVZmZmVVVVVVVVREREVVVVREREREREREREVVVVZmZmZmZmVVVVZmZmVVVVZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3d3d3ZmZmd3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3iIiIZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3d3d3d3d3ZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmiIiId3d3ZmZmd3d3VVVVREREMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREMzMzREREMzMzMzMzREREREREREREREREREREREREREREVVVVREREREREREREREREREREREREREREMzMzREREMzMzREREREREVVVVREREVVVVREREREREREREREREREREREREREREREREMzMzMzMzREREMzMzREREMzMzREREVVVVREREVVVVVVVVREREVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVREREMzMzMzMzMzMzVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmd3d3ZmZmZmZmZmZmVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREVVVVVVVVd3d3mZmZqqqqmZmZiIiId3d3d3d3VVVVREREREREVVVVVVVVVVVVd3d3ZmZmZmZmZmZmZmZmd3d3ZmZmZmZmVVVVVVVVREREVVVVVVVVZmZmVVVVVVVVREREVVVVVVVVVVVVREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzMzMzMzMzIiIiIiIiREREREREMzMzMzMzREREVVVVVVVVREREREREMzMzMzMzREREREREREREREREREREVVVVVVVVVVVVVVVVREREREREREREZmZmd3d3VVVVVVVVZmZmZmZmVVVVREREREREREREVVVVREREMzMzVVVVVVVVZmZmZmZmREREd3d3iIiIVVVVVVVVREREREREREREREREREREREREREREREREREREREREREREVVVVREREVVVVREREZmZmd3d3d3d3ZmZmVVVVZmZmVVVVVVVVZmZmiIiId3d3VVVVZmZmVVVVVVVVVVVVVVVVREREZmZmiIiId3d3d3d3d3d3VVVVREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVREREVVVVVVVVREREREREREREREREREREREREVVVVREREREREREREZmZmZmZmZmZmVVVVZmZmd3d3ZmZmZmZmVVVVVVVVREREREREVVVVVVVVZmZmVVVVVVVVVVVVREREVVVVVVVVd3d3d3d3d3d3mZmZmZmZd3d3VVVVREREVVVVZmZmZmZmZmZmZmZmd3d3d3d3iIiIqqqqzMzMu7u7qqqqqqqqqqqqu7u7mZmZiIiIiIiImZmZmZmZiIiIiIiId3d3ZmZmZmZmZmZmZmZmd3d3d3d3ZmZmVVVVZmZmiIiIqqqqmZmZiIiIiIiIiIiIiIiImZmZqqqqqqqqqqqqmZmZd3d3ZmZmZmZmVVVVZmZmVVVVVVVVZmZmZmZmd3d3iIiIiIiImZmZmZmZmZmZmZmZqqqqqqqqmZmZmZmZqqqqqqqqu7u7zMzM7u7u////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7t3d3d3d3czMzN3d3d3d3czMzMzMzN3d3czMzMzMzMzMzMzMzMzMzMzMzLu7u8zMzMzMzLu7u8zMzMzMzMzMzMzMzMzMzMzMzMzMzN3d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzLu7u7u7u6qqqpmZmaqqqqqqqqqqqqqqqqqqqru7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqru7u7u7u7u7u8zMzLu7u6qqqqqqqpmZmZmZmYiIiIiIiHd3d3d3d2ZmZmZmZlVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVURERERERDMzM0RERERERERERERERDMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERERERDMzM0RERERERERERERERERERERERFVVVVVVVVVVVWZmZmZmZlVVVWZmZmZmZlVVVVVVVVVVVXd3d2ZmZlVVVVVVVURERFVVVURERERERERERERERERERERERFVVVURERERERFVVVVVVVVVVVVVVVXd3d2ZmZlVVVVVVVWZmZmZmZmZmZmZmZnd3d2ZmZnd3d4iIiJmZmYiIiHd3d4iIiJmZmYiIiGZmZmZmZnd3d3d3d4iIiIiIiIiIiHd3d3d3d5mZmZmZmZmZmZmZmaqqqqqqqoiIiGZmZnd3d4iIiIiIiIiIiIiIiGZmZlVVVYiIiJmZmaqqqqqqqpmZmWZmZoiIiMzMzMzMzMzMzMzMzMzMzKqqqoiIiKqqqqqqqqqqqpmZmZmZmZmZmYiIiIiIiJmZmZmZmYiIiJmZmZmZmZmZmZmZmZmZmXd3d1VVVVVVVURERFVVVYiIiIiIiIiIiGZmZmZmZlVVVWZmZnd3d3d3d4iIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZnd3d4iIiIiIiHd3d3d3d4iIiHd3d4iIiIiIiHd3d4iIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiHd3d2ZmZnd3d4iIiHd3d2ZmZmZmZmZmZnd3d4iIiHd3d3d3d4iIiIiIiIiIiJmZmXd3d2ZmZlVVVVVVVWZmZnd3d3d3d2ZmZmZmZnd3d2ZmZnd3d3d3d2ZmZoiIiJmZmZmZmYiIiIiIiHd3d2ZmZmZmZmZmZnd3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d5mZmYiIiIiIiHd3d2ZmZmZmZlVVVWZmZlVVVVVVVWZmZlVVVWZmZlVVVWZmZlVVVWZmZnd3d5mZmZmZmZmZmYiIiIiIiHd3d3d3d3d3d2ZmZnd3d3d3d2ZmZlVVVWZmZlVVVVVVVWZmZoiIiIiIiHd3d3d3d3d3d3d3d1VVVWZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVURERFVVVVVVVWZmZoiIiIiIiIiIiHd3d3d3d2ZmZmZmZlVVVVVVVXd3d2ZmZlVVVVVVVWZmZmZmZlVVVVVVVXd3d3d3d4iIiIiIiIiIiIiIiIiIiGZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiHd3d3d3d3d3d2ZmZmZmZlVVVWZmZmZmZnd3d3d3d1VVVWZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d2ZmZmZmZnd3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVWZmZlVVVVVVVVVVVURERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVVVVVWZmZnd3d2ZmZlVVVWZmZlVVVVVVVVVVVWZmZlVVVVVVVURERFVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZnd3d2ZmZnd3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZlVVVWZmZlVVVWZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZnd3d2ZmZnd3d5mZmXd3d2ZmZmZmZmZmZmZmZmZmZlVVVVVVVURERFVVVVVVVVVVVVVVVVVVVURERERERFVVVURERFVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZlVVVVVVVVVVVURERERERERERERERERERERERERERERERERERDMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERDMzM0RERDMzMzMzM0RERERERERERERERERERERERERERERERERERDMzM0RERDMzM0RERERERERERERERERERERERERERFVVVURERFVVVVVVVVVVVURERFVVVURERFVVVURERERERDMzM0RERDMzM0RERERERDMzM0RERFVVVVVVVVVVVURERFVVVURERERERDMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzM0RERERERCIiIiIiIjMzM0RERFVVVVVVVVVVVWZmZlVVVWZmZmZmZnd3d2ZmZmZmZnd3d2ZmZnd3d2ZmZmZmZnd3d3d3d2ZmZmZmZlVVVURERERERERERDMzMzMzMzMzMzMzM1VVVURERERERFVVVWZmZnd3d7u7u6qqqoiIiIiIiHd3d2ZmZkRERERERFVVVVVVVWZmZnd3d2ZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZlVVVVVVVURERERERFVVVVVVVVVVVURERERERERERFVVVURERDMzM0RERERERDMzMzMzMzMzM0RERERERDMzMzMzMzMzMzMzM0RERERERDMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERFVVVVVVVURERERERERERDMzM0RERERERERERDMzM0RERERERFVVVVVVVVVVVURERERERFVVVXd3d2ZmZlVVVVVVVWZmZlVVVVVVVURERDMzMzMzM0RERDMzM0RERERERFVVVWZmZnd3d1VVVWZmZoiIiGZmZlVVVVVVVURERERERERERERERERERERERERERERERDMzM0RERERERFVVVVVVVWZmZnd3d4iIiHd3d2ZmZmZmZmZmZnd3d2ZmZlVVVVVVVWZmZnd3d3d3d3d3d2ZmZlVVVWZmZlVVVWZmZnd3d2ZmZmZmZoiIiGZmZkRERDMzM0RERERERERERFVVVVVVVURERERERFVVVURERERERERERERERFVVVXd3d3d3d1VVVVVVVVVVVURERDMzM0RERERERFVVVURERERERERERERERFVVVWZmZlVVVVVVVWZmZnd3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVURERFVVVWZmZlVVVWZmZoiIiJmZmWZmZkRERFVVVWZmZnd3d3d3d2ZmZlVVVWZmZnd3d4iIiKqqqqqqqru7u6qqqqqqqru7u6qqqqqqqqqqqpmZmXd3d4iIiIiIiIiIiHd3d3d3d3d3d2ZmZnd3d4iIiHd3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiJmZmaqqqqqqqru7u6qqqpmZmYiIiHd3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZnd3d3d3d4iIiIiIiIiIiJmZmbu7u6qqqoiIiIiIiKqqqqqqqszMzO7u7v///////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3MzMzMzMy7u7u7u7vMzMzMzMy7u7u7u7uqqqqqqqq7u7vMzMzMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7u7u7d3d3d3d3u7u7d3d3u7u7d3d3u7u7d3d3d3d3d3d3d3d3MzMzd3d3MzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7uqqqq7u7u7u7u7u7u7u7u7u7uqqqqqqqqqqqqZmZmZmZmIiIiZmZmZmZmZmZmqqqqqqqqZmZmZmZmZmZmIiIhmZmZmZmZmZmZVVVVEREREREREREQzMzNEREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzNEREQzMzNEREREREREREREREQzMzNEREREREQzMzNERERERERVVVVEREREREREREREREQzMzNEREREREREREREREREREREREREREQzMzNERERERERERERVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZmZmZmZmZVVVVmZmZVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZ3d3dVVVVVVVVmZmZ3d3d3d3d3d3d3d3dmZmZmZmZ3d3eZmZmIiIh3d3eIiIiZmZmqqqqIiIh3d3eIiIiIiIiZmZmZmZmIiIhVVVWIiIiqqqqqqqqqqqqZmZmIiIhVVVV3d3fMzMzMzMzMzMzd3d27u7uqqqqZmZmqqqqqqqq7u7u7u7uqqqqZmZmZmZmZmZl3d3eIiIiIiIiZmZmIiIiIiIiIiIiIiIh3d3dERERERERERERVVVV3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIiZmZmZmZl3d3dmZmZmZmZmZmZmZmaIiIiIiIh3d3dmZmZ3d3d3d3eIiIiIiIiIiIiIiIiZmZmqqqqZmZmIiIiIiIh3d3d3d3d3d3dmZmZmZmZ3d3dmZmZmZmZmZmZ3d3eIiIhmZmZ3d3d3d3eIiIiIiIiZmZmZmZmIiIhmZmZVVVVERERVVVVVVVVmZmZ3d3dmZmZmZmZ3d3d3d3dmZmZ3d3eZmZmZmZmIiIh3d3eIiIh3d3eIiIh3d3dVVVVmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZ3d3d3d3eIiIiZmZmIiIh3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZmZmZmZmaIiIiZmZmZmZmIiIh3d3eIiIh3d3dmZmZ3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3eIiIiIiIh3d3dmZmZmZmZVVVVVVVVVVVVVVVVmZmZVVVVmZmZVVVVERERVVVVERERVVVVmZmZ3d3eIiIiIiIh3d3d3d3dVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZVVVVmZmZVVVVVVVVmZmZmZmZ3d3eIiIiIiIh3d3eIiIh3d3dmZmZmZmZVVVVmZmZmZmZ3d3dmZmZmZmZmZmZVVVVVVVVmZmZmZmZ3d3eIiIh3d3d3d3d3d3d3d3eIiIh3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZVVVV3d3dmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVERERERERERERVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVERERVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVV3d3dmZmZVVVVVVVVERERERERERERVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3dmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmaIiIiIiIh3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVERERVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREQzMzNEREQzMzNEREQzMzNERERERERERERERERERERERERVVVVVVVVVVVVVVVVEREREREREREREREREREQzMzNEREQzMzMzMzNERERERERVVVVERERVVVVVVVVVVVVEREREREREREQzMzNEREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNERERERERVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVmZmZmZmZ3d3d3d3d3d3dmZmZVVVVEREREREQzMzMzMzNEREREREREREQzMzNERERERERmZmZ3d3eqqqq7u7uZmZmZmZmIiIh3d3dVVVVVVVVVVVVmZmZ3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVERERERERERERERERERERERERERERmZmZEREREREQzMzNERERERERERERERERERERVVVVEREQzMzMzMzMzMzMzMzNERERVVVVEREREREQzMzNEREREREREREQzMzMzMzNERERERERVVVVEREREREQzMzMzMzNEREQzMzNERERERERERERVVVVVVVVERERERERERERVVVVERERVVVVmZmZERERVVVVVVVVVVVVVVVVEREREREREREQzMzNERERERERmZmZmZmZ3d3dmZmZVVVV3d3eIiIhmZmZVVVVEREREREREREREREREREREREREREREREQzMzMzMzNERERERERERERVVVVmZmaIiIiZmZmIiIh3d3dmZmZ3d3d3d3dmZmZVVVVERERVVVV3d3eZmZmZmZl3d3dmZmZmZmZmZmZVVVV3d3eIiIhmZmaIiIh3d3dVVVVEREQzMzNERERERERERERVVVVERERVVVVERERERERVVVVERERVVVVVVVV3d3eIiIhmZmZVVVVVVVVERERERERERERERERERERERERERERmZmZVVVVVVVVVVVVVVVVERERVVVV3d3d3d3dVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVERERmZmaIiIhVVVVmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmaIiIiqqqq7u7uqqqqqqqq7u7vMzMy7u7uqqqqqqqqZmZl3d3d3d3eZmZmqqqqIiIiZmZmZmZmqqqqZmZmZmZmqqqqqqqqqqqqZmZmZmZmZmZmZmZmqqqqqqqqqqqqqqqqZmZmIiIhmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVmZmZVVVVVVVV3d3eIiIiIiIiZmZmqqqqZmZmIiIh3d3eZmZm7u7vMzMzd3d3///////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3dzMzM3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMu7u7zMzMzMzMzMzMzMzMzMzM3d3d3d3d3d3d7u7u7u7u3d3d7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7zMzMu7u7u7u7u7u7qqqqu7u7u7u7qqqqmZmZiIiId3d3ZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmVVVVVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREREREREREREREMzMzREREMzMzREREREREREREMzMzREREMzMzMzMzMzMzREREMzMzREREMzMzREREMzMzREREREREMzMzREREMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzREREREREREREREREREREREREVVVVREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3ZmZmd3d3d3d3ZmZmVVVVVVVVZmZmVVVVREREVVVVVVVVVVVVVVVVREREREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVd3d3ZmZmZmZmZmZmZmZmZmZmZmZmiIiId3d3VVVVZmZmiIiIiIiImZmZiIiId3d3d3d3d3d3iIiImZmZZmZmZmZmqqqqmZmZmZmZqqqqmZmZZmZmREREd3d3qqqqqqqqzMzMzMzMzMzMu7u7u7u7zMzMu7u7zMzMzMzMu7u7u7u7u7u7mZmZd3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiId3d3VVVVREREVVVVZmZmd3d3ZmZmZmZmd3d3iIiId3d3d3d3d3d3d3d3iIiId3d3iIiImZmZmZmZqqqqu7u7qqqqiIiId3d3ZmZmZmZmZmZmZmZmiIiId3d3ZmZmd3d3d3d3iIiIiIiImZmZmZmZmZmZmZmZmZmZiIiId3d3d3d3d3d3iIiIZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3iIiId3d3iIiIiIiImZmZd3d3d3d3ZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVZmZmZmZmd3d3mZmZmZmZiIiIiIiIiIiIiIiIiIiIiIiIVVVVVVVVZmZmd3d3ZmZmd3d3ZmZmZmZmd3d3d3d3d3d3mZmZiIiIiIiId3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3iIiImZmZiIiIiIiIiIiId3d3d3d3ZmZmd3d3ZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3ZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVREREVVVVd3d3iIiIiIiId3d3d3d3ZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmVVVVVVVVZmZmd3d3iIiIiIiId3d3d3d3d3d3iIiId3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmiIiId3d3d3d3ZmZmZmZmVVVVZmZmZmZmVVVVZmZmZmZmd3d3d3d3ZmZmVVVVZmZmZmZmd3d3ZmZmVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREREREVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmZmZmVVVVVVVVREREVVVVREREVVVVVVVVZmZmZmZmVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREZmZmZmZmZmZmZmZmREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3ZmZmd3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmiIiIiIiIZmZmd3d3ZmZmd3d3ZmZmd3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3ZmZmd3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmd3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmVVVVZmZmVVVVZmZmZmZmVVVVVVVVVVVVZmZmZmZmd3d3ZmZmd3d3ZmZmd3d3d3d3iIiIiIiId3d3ZmZmVVVVREREMzMzREREREREMzMzREREMzMzMzMzREREREREREREVVVVVVVVVVVVREREMzMzMzMzREREMzMzREREMzMzREREREREMzMzMzMzREREMzMzREREMzMzREREMzMzREREMzMzREREREREVVVVVVVVVVVVREREREREREREVVVVREREREREREREMzMzREREMzMzMzMzREREREREVVVVVVVVVVVVVVVVVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzREREREREVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREMzMzMzMzMzMzREREREREZmZmiIiIu7u7qqqqqqqqmZmZiIiIZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmd3d3ZmZmZmZmZmZmZmZmVVVVVVVVREREREREREREREREREREVVVVZmZmREREREREMzMzREREREREREREVVVVREREREREREREMzMzREREREREREREREREVVVVREREREREMzMzMzMzREREREREREREIiIiMzMzREREREREREREREREREREMzMzMzMzMzMzIiIiMzMzVVVVVVVVREREREREREREVVVVREREREREVVVVVVVVVVVVVVVVVVVVREREREREREREMzMzREREREREVVVVVVVVVVVVVVVVZmZmVVVVREREiIiIiIiIZmZmVVVVVVVVVVVVREREREREREREREREREREREREMzMzREREMzMzREREREREZmZmVVVVd3d3mZmZiIiIZmZmZmZmd3d3ZmZmVVVVREREREREREREZmZmd3d3iIiIiIiIZmZmZmZmZmZmZmZmiIiImZmZZmZmiIiIiIiIZmZmREREMzMzREREMzMzREREREREREREREREVVVVVVVVREREVVVVVVVVVVVVVVVVd3d3d3d3ZmZmVVVVREREMzMzREREREREREREREREREREVVVVVVVVREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVd3d3ZmZmd3d3VVVVVVVVREREREREVVVVVVVVVVVVVVVVZmZmiIiIVVVVVVVVZmZmZmZmZmZmiIiId3d3ZmZmZmZmZmZmd3d3d3d3d3d3d3d3mZmZqqqqqqqqu7u73d3d3d3dzMzMqqqqmZmZiIiId3d3iIiIqqqqqqqqqqqqmZmZqqqqu7u7mZmZmZmZu7u7qqqqmZmZmZmZmZmZiIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmZmZmd3d3ZmZmZmZmVVVVZmZmZmZmVVVVZmZmVVVVVVVVZmZmVVVVZmZmZmZmd3d3mZmZmZmZiIiId3d3d3d3mZmZu7u7zMzM3d3d7u7u////////7u7u////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7t3d3d3d3d3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzLu7u8zMzLu7u7u7u6qqqpmZmaqqqpmZmZmZmYiIiHd3d2ZmZlVVVURERERERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMzMzM0RERERERDMzM0RERDMzM0RERERERERERFVVVURERERERERERERERERERERERERERDMzM0RERERERERERDMzM0RERDMzMzMzM0RERERERDMzM0RERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVXd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVURERERERERERERERERERFVVVWZmZmZmZnd3d3d3d2ZmZnd3d4iIiHd3d2ZmZlVVVWZmZmZmZnd3d3d3d3d3d5mZmWZmZlVVVVVVVWZmZmZmZoiIiJmZmWZmZmZmZmZmZoiIiHd3d1VVVXd3d6qqqpmZmZmZmaqqqpmZmXd3d1VVVXd3d6qqqqqqqru7u93d3czMzLu7u8zMzMzMzLu7u7u7u93d3czMzLu7u7u7u5mZmXd3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d2ZmZnd3d3d3d3d3d2ZmZmZmZlVVVWZmZoiIiIiIiHd3d2ZmZnd3d3d3d3d3d3d3d5mZmZmZmZmZmZmZmaqqqpmZmZmZmYiIiHd3d2ZmZmZmZnd3d3d3d3d3d3d3d2ZmZnd3d4iIiIiIiKqqqpmZmZmZmaqqqnd3d3d3d4iIiIiIiIiIiIiIiFVVVWZmZmZmZnd3d3d3d4iIiHd3d2ZmZoiIiIiIiIiIiHd3d4iIiJmZmXd3d3d3d2ZmZlVVVURERFVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZpmZmZmZmYiIiHd3d3d3d4iIiIiIiHd3d2ZmZlVVVWZmZlVVVWZmZmZmZnd3d2ZmZnd3d2ZmZoiIiIiIiIiIiHd3d3d3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZlVVVURERFVVVWZmZmZmZmZmZoiIiIiIiHd3d4iIiHd3d3d3d2ZmZmZmZnd3d2ZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZmZmZnd3d3d3d3d3d3d3d3d3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVWZmZmZmZnd3d4iIiHd3d4iIiHd3d3d3d4iIiIiIiHd3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d4iIiGZmZlVVVWZmZlVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZlVVVVVVVVVVVXd3d3d3d2ZmZlVVVVVVVVVVVURERFVVVURERFVVVVVVVURERFVVVWZmZmZmZmZmZlVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVURERFVVVURERERERGZmZlVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVXd3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVVVVVWZmZmZmZlVVVVVVVVVVVURERFVVVVVVVVVVVURERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d3d3d3d3d2ZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZnd3d2ZmZmZmZnd3d2ZmZnd3d2ZmZnd3d4iIiHd3d2ZmZmZmZnd3d2ZmZnd3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZoiIiIiIiHd3d3d3d3d3d3d3d2ZmZnd3d2ZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZlVVVVVVVWZmZlVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d2ZmZnd3d2ZmZnd3d2ZmZmZmZnd3d2ZmZnd3d2ZmZnd3d2ZmZmZmZmZmZlVVVWZmZlVVVWZmZlVVVWZmZmZmZlVVVWZmZmZmZnd3d2ZmZnd3d3d3d4iIiHd3d2ZmZlVVVWZmZmZmZmZmZmZmZlVVVVVVVURERDMzM0RERERERFVVVURERERERERERERERDMzM0RERERERERERERERDMzM0RERDMzMzMzMzMzMzMzM0RERERERDMzM0RERDMzM0RERDMzM1VVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERDMzMzMzM0RERFVVVURERFVVVVVVVVVVVURERERERDMzMzMzM0RERERERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVVVVVVVVVVVVVWZmZnd3d2ZmZmZmZlVVVWZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZlVVVURERERERDMzMzMzMzMzM1VVVVVVVYiIiLu7u7u7u6qqqpmZmYiIiHd3d1VVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVWZmZnd3d2ZmZnd3d2ZmZmZmZkRERERERERERERERDMzM0RERFVVVURERERERDMzM0RERERERERERFVVVURERERERERERERERDMzM0RERFVVVURERERERERERERERERERDMzMzMzMzMzM0RERERERDMzMzMzM0RERERERERERERERDMzMzMzM0RERDMzMzMzMzMzM0RERGZmZlVVVURERERERERERERERDMzM0RERFVVVURERFVVVURERFVVVVVVVURERDMzMzMzM1VVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVYiIiJmZmWZmZlVVVVVVVURERERERERERERERERERERERDMzM0RERERERERERERERERERFVVVVVVVXd3d4iIiIiIiGZmZlVVVWZmZmZmZlVVVVVVVURERFVVVURERGZmZmZmZmZmZmZmZlVVVVVVVWZmZoiIiJmZmXd3d3d3d4iIiGZmZkRERDMzM0RERERERDMzM0RERERERFVVVVVVVVVVVURERFVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZkRERDMzM0RERERERERERERERERERDMzM0RERDMzM0RERERERERERERERFVVVVVVVVVVVVVVVVVVVXd3d3d3d3d3d1VVVVVVVVVVVURERFVVVURERFVVVWZmZnd3d5mZmWZmZmZmZnd3d2ZmZnd3d3d3d3d3d2ZmZlVVVWZmZoiIiGZmZnd3d4iIiIiIiIiIiKqqqru7u7u7u93d3d3d3aqqqoiIiIiIiHd3d5mZmaqqqru7u6qqqoiIiJmZmaqqqpmZmYiIiIiIiHd3d3d3d4iIiHd3d4iIiHd3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZnd3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVXd3d4iIiIiIiHd3d3d3d3d3d4iIiKqqqru7u8zMzO7u7v///////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7u7u7d3d3d3d3u7u7d3d3u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3MzMzMzMy7u7u7u7u7u7uZmZmIiIiIiIh3d3d3d3dmZmZVVVVVVVVEREREREQzMzMzMzNEREQzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNEREREREREREQzMzMzMzNERERVVVVERERERERERERERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVERERVVVVEREREREQzMzMzMzNERERVVVVmZmaIiIh3d3d3d3eIiIiIiIh3d3d3d3eIiIiIiIh3d3dVVVVVVVVmZmZ3d3eIiIiIiIiIiIhmZmZVVVVVVVVVVVVmZmZ3d3d3d3dVVVVVVVVmZmZmZmZVVVVVVVWZmZmqqqqZmZmqqqqqqqqIiIiIiIhmZmZmZmaqqqq7u7vMzMzMzMzMzMy7u7vMzMzMzMy7u7vMzMzMzMzMzMy7u7u7u7uZmZmIiIiIiIhmZmZmZmZmZmZmZmZmZmZ3d3d3d3eIiIiZmZmZmZmIiIhmZmZ3d3dmZmZmZmaIiIh3d3dmZmZ3d3d3d3d3d3eIiIiZmZmqqqqIiIiIiIiZmZmIiIiIiIh3d3dmZmZmZmZmZmZ3d3d3d3d3d3d3d3dmZmZ3d3d3d3eZmZmqqqqqqqqZmZmIiIh3d3d3d3eIiIiZmZmZmZmIiIhmZmZmZmZ3d3d3d3eIiIiIiIh3d3d3d3d3d3eIiIh3d3eIiIiIiIiIiIh3d3d3d3dmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZVVVVmZmZmZmZmZmZ3d3d3d3d3d3eIiIiIiIiIiIh3d3dmZmZmZmZmZmZVVVVmZmZVVVVVVVVmZmZ3d3dmZmZVVVVERERVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3dmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZmZmaIiIh3d3d3d3dmZmZ3d3d3d3dmZmZVVVVVVVVVVVVmZmZmZmZVVVVVVVVmZmZmZmZ3d3dmZmZmZmZmZmZVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVmZmaIiIiIiIh3d3dmZmZmZmZmZmZ3d3eIiIiIiIhmZmZmZmZVVVVVVVVVVVVERERVVVVmZmZVVVVVVVVmZmZVVVVmZmZVVVVmZmZmZmZmZmZmZmZ3d3dVVVVmZmZVVVVmZmZmZmZmZmZVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZVVVVVVVVmZmZ3d3d3d3dVVVVERERERERVVVVERERERERVVVVVVVVERERERERERERmZmZ3d3dmZmZVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVERERVVVVERERVVVVVVVVmZmZVVVVVVVVVVVVEREQzMzNERERERERERERERERVVVVVVVVmZmZVVVVmZmZVVVVmZmZVVVV3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVERERVVVVERERVVVVVVVVERERERERVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZ3d3dmZmZ3d3d3d3dmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZ3d3eIiIiIiIh3d3eIiIh3d3d3d3d3d3eIiIh3d3d3d3d3d3d3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZ3d3d3d3dmZmZ3d3dmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3eIiIh3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZ3d3d3d3dmZmZ3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZ3d3dmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3dmZmZmZmZmZmZmZmZVVVVEREREREQzMzNEREQzMzMzMzNEREQzMzMzMzNEREQzMzNEREQzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzNERERERERVVVVVVVVVVVVVVVVVVVVEREQzMzNEREREREREREREREQzMzNEREQzMzNERERVVVVERERERERVVVVVVVVVVVVEREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVVVVVVVVVVVVVmZmZ3d3d3d3dmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZVVVV3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVUzMzMzMzMzMzMzMzNERERVVVV3d3eqqqq7u7uqqqqZmZmZmZmZmZl3d3dVVVVmZmZmZmZVVVVVVVVERERVVVVVVVVmZmZmZmZmZmZmZmZ3d3dmZmZEREREREQzMzMzMzNERERERERVVVVEREQzMzNERERERERERERERERVVVVEREREREREREREREREREQzMzNERERERERERERERERVVVVEREQzMzMzMzMzMzNEREREREQzMzMzMzMzMzNEREREREREREREREQzMzMzMzNEREQzMzMzMzNERERVVVVEREREREQzMzNEREQzMzNERERERERERERVVVVVVVVERERERERVVVUzMzMzMzMzMzNERERmZmZmZmZVVVVmZmZVVVVVVVVVVVV3d3eIiIhmZmZVVVVVVVVEREREREREREREREQzMzNEREQzMzMzMzNERERERERERERERERVVVVVVVVmZmZ3d3eIiIhmZmZVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERmZmZVVVVmZmZmZmZ3d3eIiIiIiIiIiIiIiIiIiIhmZmZEREREREQzMzNERERERERERERERERVVVVmZmZVVVVVVVVERERERERERERERERERERERERmZmZmZmZVVVUzMzNEREQzMzNEREQzMzNEREREREQzMzNERERERERERERERERERERERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVERERERERVVVVVVVVmZmZ3d3dmZmZ3d3eIiIh3d3eIiIiIiIhmZmZ3d3dmZmZmZmZ3d3eIiIh3d3eIiIh3d3d3d3e7u7u7u7uqqqq7u7u7u7uIiIiIiIiqqqqZmZmZmZmqqqrMzMy7u7uIiIiIiIiZmZmIiIiIiIh3d3d3d3dmZmZ3d3d3d3eIiIh3d3d3d3eIiIh3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZ3d3d3d3dVVVVmZmZmZmZ3d3d3d3eIiIiIiIiIiIiqqqq7u7vMzMzd3d3///////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d7u7u3d3d7u7u7u7u3d3d7u7u3d3d7u7u3d3d7u7u3d3d7u7u3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3du7u7mZmZiIiIiIiId3d3VVVVVVVVREREREREREREMzMzMzMzMzMzREREREREREREREREREREREREREREVVVVREREREREVVVVREREREREVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmd3d3ZmZmZmZmd3d3ZmZmd3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3iIiIiIiIiIiImZmZmZmZiIiIiIiImZmZiIiIiIiIiIiId3d3d3d3d3d3d3d3ZmZmd3d3ZmZmZmZmd3d3d3d3ZmZmVVVVZmZmZmZmd3d3d3d3ZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREREREREREREREREREVVVVREREREREREREREREMzMzREREMzMzMzMzREREMzMzMzMzMzMzMzMzVVVVd3d3d3d3iIiIiIiIiIiIZmZmVVVVd3d3d3d3d3d3d3d3iIiIZmZmZmZmVVVVZmZmZmZmiIiId3d3ZmZmZmZmd3d3d3d3ZmZmVVVVVVVVZmZmZmZmVVVVZmZmZmZmZmZmd3d3qqqqzMzMu7u7qqqqqqqqd3d3d3d3ZmZmd3d3mZmZzMzM3d3dzMzMu7u7u7u7zMzMu7u7u7u7u7u7u7u7qqqqmZmZmZmZmZmZmZmZiIiId3d3ZmZmREREVVVVVVVVd3d3mZmZmZmZmZmZd3d3iIiId3d3ZmZmd3d3d3d3d3d3ZmZmZmZmd3d3ZmZmd3d3mZmZqqqqqqqqmZmZiIiIiIiIiIiIiIiId3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3iIiId3d3iIiImZmZqqqqmZmZmZmZiIiId3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3iIiId3d3d3d3iIiId3d3d3d3d3d3d3d3iIiId3d3iIiIiIiId3d3d3d3VVVVZmZmd3d3ZmZmZmZmZmZmiIiIiIiId3d3d3d3d3d3iIiIiIiId3d3d3d3ZmZmZmZmZmZmZmZmd3d3ZmZmVVVVVVVVVVVVZmZmZmZmd3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmVVVVVVVVZmZmZmZmVVVVVVVVZmZmVVVVVVVVREREVVVVZmZmZmZmZmZmd3d3d3d3iIiId3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmVVVVZmZmZmZmd3d3d3d3d3d3d3d3d3d3iIiId3d3ZmZmZmZmZmZmVVVVVVVVZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVREREVVVVREREVVVVREREVVVVREREVVVVVVVVZmZmVVVVVVVVREREREREVVVVZmZmd3d3d3d3ZmZmVVVVVVVVVVVVZmZmd3d3d3d3d3d3ZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmd3d3iIiIZmZmZmZmZmZmVVVVZmZmVVVVREREVVVVREREVVVVZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmVVVVVVVVREREVVVVREREREREREREVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVREREREREREREVVVVVVVVVVVVZmZmVVVVVVVVREREREREREREREREREREVVVVREREVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmd3d3ZmZmZmZmVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVd3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmVVVVZmZmZmZmVVVVZmZmVVVVZmZmZmZmd3d3d3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmVVVVZmZmVVVVZmZmVVVVZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiId3d3iIiIiIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmd3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmd3d3d3d3d3d3d3d3iIiIiIiIiIiId3d3iIiIiIiIiIiId3d3ZmZmZmZmVVVVVVVVREREREREMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVVVVVVVVVVVVVREREREREREREREREREREMzMzREREMzMzMzMzMzMzREREREREREREVVVVVVVVVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREVVVVVVVVVVVVZmZmd3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVd3d3d3d3ZmZmZmZmVVVVZmZmZmZmZmZmVVVVVVVVREREREREVVVVMzMzMzMzREREVVVVZmZmiIiIu7u7qqqqqqqqqqqqqqqqiIiId3d3d3d3ZmZmVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3ZmZmVVVVMzMzMzMzMzMzMzMzVVVVVVVVVVVVREREMzMzREREMzMzMzMzREREVVVVVVVVREREVVVVREREVVVVREREREREREREVVVVVVVVREREMzMzREREMzMzREREREREMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzREREMzMzMzMzREREREREVVVVVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzVVVVZmZmZmZmVVVVZmZmVVVVREREREREd3d3mZmZZmZmZmZmVVVVREREREREREREREREREREMzMzREREREREREREREREREREREREREREREREZmZmd3d3ZmZmVVVVVVVVZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmd3d3iIiIiIiId3d3mZmZmZmZVVVVREREREREREREREREREREVVVVVVVVREREVVVVZmZmREREVVVVREREREREREREREREREREVVVVVVVVVVVVMzMzMzMzREREMzMzREREREREMzMzREREREREMzMzREREREREREREREREVVVVVVVVZmZmVVVVREREREREREREZmZmd3d3ZmZmVVVVZmZmZmZmVVVVVVVVREREVVVVZmZmd3d3d3d3d3d3iIiIiIiIiIiId3d3d3d3ZmZmd3d3iIiId3d3d3d3ZmZmd3d3mZmZmZmZmZmZqqqqiIiIiIiImZmZu7u7zMzMqqqqu7u7zMzMu7u7u7u7u7u7mZmZiIiId3d3d3d3d3d3d3d3iIiIiIiId3d3d3d3iIiIiIiId3d3ZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3iIiImZmZqqqqu7u73d3d3d3d////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////+7u7v///////+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7t3d3e7u7t3d3e7u7t3d3e7u7u7u7t3d3e7u7t3d3d3d3d3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3czMzLu7u7u7u5mZmYiIiGZmZlVVVVVVVURERERERERERERERERERERERERERFVVVVVVVVVVVWZmZmZmZmZmZnd3d2ZmZnd3d3d3d3d3d2ZmZnd3d2ZmZlVVVXd3d2ZmZnd3d3d3d3d3d3d3d4iIiHd3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d4iIiHd3d4iIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiIiIiIiIiHd3d3d3d2ZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMyIiIjMzMyIiIiIiIjMzMzMzM0RERFVVVXd3d3d3d4iIiIiIiGZmZlVVVVVVVURERGZmZmZmZnd3d3d3d3d3d3d3d2ZmZnd3d2ZmZmZmZmZmZmZmZnd3d3d3d4iIiIiIiGZmZmZmZlVVVXd3d2ZmZmZmZpmZmYiIiIiIiLu7u8zMzLu7u7u7u7u7u3d3d2ZmZnd3d4iIiJmZmczMzMzMzMzMzJmZmbu7u7u7u6qqqqqqqqqqqqqqqqqqqpmZmaqqqpmZmYiIiIiIiIiIiHd3d3d3d2ZmZlVVVXd3d6qqqpmZmZmZmYiIiIiIiHd3d2ZmZnd3d4iIiGZmZmZmZmZmZmZmZmZmZnd3d4iIiJmZmZmZmYiIiIiIiHd3d4iIiHd3d3d3d3d3d2ZmZnd3d3d3d3d3d2ZmZnd3d4iIiIiIiJmZmZmZmZmZmZmZmYiIiIiIiHd3d4iIiHd3d3d3d4iIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiHd3d5mZmZmZmYiIiHd3d3d3d2ZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d2ZmZlVVVVVVVWZmZlVVVVVVVWZmZmZmZnd3d3d3d2ZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZlVVVURERFVVVVVVVVVVVWZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZlVVVURERFVVVWZmZnd3d2ZmZmZmZnd3d4iIiHd3d3d3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVURERFVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVURERFVVVWZmZmZmZnd3d2ZmZlVVVWZmZlVVVWZmZmZmZnd3d3d3d1VVVWZmZlVVVWZmZkRERFVVVURERERERGZmZmZmZmZmZmZmZlVVVVVVVWZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVURERERERDMzM0RERFVVVWZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVURERFVVVURERERERERERFVVVVVVVVVVVURERERERERERERERFVVVVVVVWZmZmZmZlVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVURERDMzM0RERERERFVVVWZmZmZmZmZmZkRERERERERERERERFVVVURERERERERERERERFVVVVVVVURERFVVVVVVVURERERERERERERERFVVVVVVVWZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVWZmZlVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d2ZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiHd3d4iIiIiIiIiIiJmZmYiIiIiIiHd3d2ZmZnd3d3d3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d2ZmZnd3d3d3d2ZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiHd3d4iIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d3d3d2ZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d4iIiJmZmYiIiIiIiIiIiIiIiHd3d4iIiIiIiHd3d2ZmZmZmZmZmZlVVVVVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVVVVVURERERERERERERERDMzM0RERDMzM0RERERERDMzMzMzMzMzM0RERERERERERERERFVVVVVVVTMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzM0RERERERERERERERFVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVVVVVWZmZmZmZnd3d2ZmZlVVVWZmZnd3d3d3d3d3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVYiIiKqqqru7u6qqqqqqqqqqqoiIiIiIiGZmZlVVVVVVVVVVVVVVVVVVVVVVVURERFVVVWZmZmZmZlVVVWZmZlVVVVVVVTMzMzMzMzMzM0RERFVVVVVVVURERERERDMzM0RERDMzMzMzM0RERERERERERERERFVVVURERERERERERERERFVVVVVVVURERERERDMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERDMzM0RERERERERERERERDMzMzMzMzMzM0RERERERFVVVVVVVURERDMzMyIiIjMzMzMzMzMzM0RERGZmZnd3d3d3d3d3d1VVVVVVVVVVVURERGZmZoiIiHd3d1VVVVVVVVVVVURERERERERERERERFVVVURERERERERERERERDMzM0RERERERFVVVWZmZmZmZmZmZmZmZlVVVVVVVVVVVXd3d3d3d3d3d3d3d4iIiHd3d3d3d4iIiHd3d2ZmZlVVVWZmZoiIiHd3d4iIiJmZmYiIiHd3d1VVVVVVVWZmZlVVVWZmZmZmZmZmZlVVVURERFVVVURERFVVVURERERERFVVVVVVVVVVVURERFVVVVVVVURERDMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERERERERERERERERERFVVVWZmZmZmZlVVVVVVVVVVVWZmZoiIiHd3d2ZmZmZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZnd3d2ZmZoiIiJmZmYiIiHd3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d4iIiJmZmZmZmXd3d3d3d3d3d5mZmczMzMzMzLu7u6qqqqqqqru7u6qqqqqqqoiIiIiIiHd3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiHd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZnd3d2ZmZmZmZmZmZmZmZnd3d3d3d4iIiIiIiIiIiJmZmaqqqqqqqqqqqszMzO7u7u7u7v///////+7u7v///////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3u7u7d3d3d3d3d3d3u7u7u7u7d3d3d3d3MzMzMzMzMzMzMzMzd3d3d3d3MzMzd3d3MzMzd3d3MzMzd3d3MzMy7u7u7u7u7u7uZmZmIiIh3d3d3d3dmZmZVVVVERERERERERERVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3eIiIh3d3eIiIiIiIiZmZmIiIh3d3eIiIiIiIiIiIh3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZVVVVmZmZVVVVVVVVmZmZVVVVmZmZmZmZ3d3eIiIh3d3d3d3d3d3eIiIh3d3d3d3dmZmZmZmZmZmZVVVVVVVVERERVVVVVVVVEREREREQzMzMzMzMzMzMiIiIiIiIiIiIzMzMiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzNERERVVVVVVVVVVVVmZmZmZmZ3d3dmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZ3d3eIiIh3d3d3d3d3d3d3d3dVVVVmZmaIiIiZmZmIiIiIiIiZmZmIiIhmZmZVVVVmZmZmZmZ3d3eIiIh3d3eIiIiqqqrd3d3MzMzMzMyqqqqIiIhVVVV3d3eIiIiIiIiqqqq7u7uqqqqqqqq7u7u7u7uZmZm7u7uqqqqqqqq7u7uqqqqqqqqqqqqIiIiIiIiIiIiIiIiIiIh3d3dVVVV3d3eZmZmZmZmZmZmIiIiIiIh3d3dmZmZ3d3d3d3d3d3dmZmZmZmZmZmZmZmaIiIiZmZmZmZmIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3dVVVVmZmZmZmZmZmZmZmZmZmZ3d3eZmZmZmZmIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3eIiIh3d3d3d3eIiIh3d3d3d3d3d3dmZmZmZmZ3d3eIiIiZmZmZmZmIiIiIiIiZmZmZmZl3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3eIiIh3d3d3d3eIiIiIiIiIiIh3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVVVVVmZmZVVVVVVVVmZmZ3d3dmZmZmZmZmZmaIiIh3d3dmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVV3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVVVVVmZmZVVVVERERERERVVVVmZmZmZmZmZmZmZmZ3d3d3d3dmZmZmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVERERVVVVVVVVERERERERVVVVVVVVVVVVVVVVERERVVVVmZmZVVVVERERERERERERVVVV3d3dmZmZVVVVmZmZmZmZ3d3dmZmZVVVVmZmZmZmZmZmZmZmZ3d3dmZmZVVVVVVVVERERERERERERVVVVVVVVmZmZmZmZmZmZmZmZ3d3d3d3d3d3dmZmZmZmZmZmZVVVVmZmZVVVVEREQzMzMzMzNERERVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVVVVVVVVVERERERERERERERERVVVVVVVVmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVERERVVVVmZmZVVVVVVVVVVVVEREREREQzMzNERERERERVVVVmZmZmZmZVVVVERERERERERERVVVUzMzNERERERERERERVVVVVVVVEREREREREREREREQzMzMzMzNERERVVVVVVVVVVVVERERVVVVmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3eZmZmZmZmIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIh3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3eIiIiIiIiZmZmIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3dmZmZ3d3dmZmZ3d3dmZmZ3d3d3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZ3d3d3d3eIiIiZmZmqqqqZmZmIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3dmZmZVVVVVVVUzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVVVVVEREREREREREREREREREREREQzMzNEREQzMzMzMzMzMzMzMzNERERERERERERERERVVVVVVVVEREREREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERVVVVVVVVVVVVmZmZmZmZ3d3dmZmZmZmZVVVVVVVVVVVVVVVVmZmZ3d3dmZmZ3d3dmZmZmZmZVVVVmZmaIiIh3d3d3d3dmZmZmZmZERERERERVVVVmZmZmZmZERERERERVVVV3d3eqqqq7u7u7u7uZmZmIiIiZmZmIiIh3d3dVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVUzMzMzMzNEREQzMzNERERVVVVEREREREREREQzMzMzMzMzMzNEREQzMzNERERVVVVERERERERERERERERERERERERVVVVEREQzMzNEREQzMzNEREQzMzNEREQzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNERERERERVVVVVVVVEREQzMzMzMzNEREQzMzMzMzNERERVVVVVVVVVVVUzMzMiIiIzMzMzMzMzMzNERERVVVWIiIiZmZl3d3dmZmZVVVVERERERERmZmaZmZl3d3d3d3dVVVVEREREREREREQzMzNEREREREREREQzMzNEREQzMzNERERERERVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVmZmZ3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIh3d3dmZmZ3d3eIiIiIiIiIiIh3d3eIiIiZmZmZmZlmZmZmZmZVVVVmZmZmZmZ3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZVVVVEREREREQzMzNEREQzMzMzMzMzMzNERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3dmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZ3d3d3d3dmZmZ3d3d3d3d3d3dmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmaIiIiIiIh3d3dmZmZmZmZ3d3eIiIiqqqqqqqqqqqqIiIiqqqqqqqqZmZmIiIh3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiZmZmIiIh3d3dmZmZVVVVVVVVVVVVmZmZ3d3eIiIiIiIhmZmZVVVVmZmZ3d3d3d3dmZmZ3d3d3d3eIiIiIiIiZmZmZmZmZmZmZmZm7u7u7u7u7u7vd3d3u7u7///////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3d3d3dzMzM3d3dzMzMu7u7qqqqqqqqqqqqqqqqu7u7u7u7u7u7u7u7zMzMzMzMzMzMzMzMu7u7zMzMzMzMu7u7qqqqiIiIiIiId3d3ZmZmd3d3ZmZmd3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiImZmZqqqqmZmZmZmZmZmZiIiIiIiIiIiId3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3iIiIiIiIiIiImZmZmZmZmZmZmZmZiIiId3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiId3d3d3d3ZmZmZmZmZmZmZmZmREREREREREREREREMzMzREREMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzIiIiIiIiMzMzIiIiMzMzMzMzREREMzMzIiIiIiIiMzMzMzMzMzMzREREZmZmZmZmVVVVVVVVZmZmZmZmZmZmVVVVZmZmZmZmZmZmiIiImZmZd3d3ZmZmd3d3mZmZd3d3ZmZmd3d3d3d3d3d3ZmZmiIiImZmZiIiIiIiImZmZiIiId3d3ZmZmZmZmZmZmiIiImZmZd3d3d3d3iIiIu7u7zMzMqqqqmZmZiIiIiIiId3d3iIiImZmZiIiIiIiIqqqqu7u7zMzMu7u7qqqqqqqqqqqqqqqqu7u7zMzMu7u7qqqqiIiId3d3ZmZmd3d3iIiId3d3d3d3qqqqmZmZiIiImZmZmZmZiIiIiIiIZmZmd3d3iIiIiIiIZmZmZmZmZmZmd3d3mZmZiIiIiIiIiIiIiIiIiIiImZmZiIiId3d3iIiIZmZmZmZmZmZmZmZmVVVVVVVVVVVVd3d3d3d3iIiIiIiId3d3VVVVZmZmZmZmd3d3iIiId3d3d3d3d3d3d3d3iIiIiIiId3d3ZmZmVVVVREREVVVVVVVVd3d3iIiImZmZiIiIiIiId3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmd3d3d3d3d3d3iIiImZmZiIiIiIiIiIiIiIiId3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmVVVVVVVVZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVREREVVVVREREREREREREVVVVVVVVd3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmZmZmZmZmZmZmVVVVVVVVREREMzMzREREVVVVZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVVVVVVVVVREREREREREREREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmVVVVREREMzMzREREVVVVZmZmVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVd3d3ZmZmZmZmVVVVVVVVREREMzMzMzMzREREVVVVVVVVVVVVZmZmVVVVZmZmd3d3d3d3ZmZmd3d3ZmZmVVVVZmZmZmZmVVVVREREREREMzMzREREVVVVVVVVZmZmZmZmVVVVVVVVVVVVREREVVVVREREVVVVREREREREVVVVVVVVVVVVREREREREREREMzMzREREREREVVVVZmZmVVVVREREVVVVVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREMzMzREREREREVVVVZmZmVVVVVVVVVVVVREREREREREREREREMzMzREREREREVVVVVVVVREREREREREREREREMzMzIiIiREREREREREREREREREREREREVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVd3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmd3d3iIiId3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiImZmZiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3iIiId3d3d3d3d3d3ZmZmd3d3ZmZmd3d3ZmZmd3d3d3d3d3d3ZmZmd3d3d3d3d3d3iIiId3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3ZmZmd3d3ZmZmd3d3ZmZmZmZmd3d3ZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmd3d3mZmZqqqqmZmZiIiIiIiIiIiIiIiIiIiIiIiImZmZiIiImZmZiIiImZmZiIiIiIiIiIiId3d3ZmZmVVVVMzMzMzMzMzMzMzMzMzMzIiIiMzMzREREREREREREVVVVREREREREREREREREREREMzMzREREMzMzMzMzMzMzMzMzREREREREVVVVREREREREREREREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVREREREREVVVVZmZmVVVVZmZmd3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVd3d3ZmZmZmZmZmZmVVVVZmZmd3d3iIiId3d3VVVVZmZmZmZmREREREREREREVVVVd3d3ZmZmVVVVVVVVVVVViIiIqqqqu7u7iIiIiIiIiIiImZmZd3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREMzMzMzMzMzMzREREVVVVREREREREMzMzREREREREMzMzMzMzMzMzMzMzREREREREREREREREMzMzREREREREREREREREREREREREVVVVREREMzMzREREREREREREMzMzMzMzMzMzIiIiIiIiMzMzMzMzREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVVVVVMzMzIiIiMzMzIiIiMzMzMzMzREREREREVVVVd3d3d3d3VVVVVVVVVVVVREREVVVVd3d3d3d3ZmZmZmZmREREREREMzMzREREMzMzREREMzMzREREMzMzMzMzMzMzREREMzMzREREVVVVVVVVREREVVVVZmZmZmZmZmZmd3d3iIiIiIiImZmZmZmZmZmZmZmZmZmZmZmZiIiIqqqqqqqqmZmZmZmZiIiIiIiIiIiIu7u7mZmZd3d3ZmZmVVVVd3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmd3d3d3d3VVVVVVVVREREREREREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmd3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmd3d3iIiIiIiIiIiIiIiImZmZmZmZiIiId3d3d3d3d3d3iIiIiIiImZmZiIiIiIiIiIiId3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmd3d3iIiId3d3ZmZmVVVVZmZmd3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiImZmZqqqqqqqqu7u7zMzM3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3e7u7t3d3e7u7u7u7t3d3e7u7u7u7t3d3d3d3czMzMzMzMzMzLu7u7u7u6qqqpmZmZmZmZmZmZmZmaqqqqqqqszMzMzMzMzMzMzMzMzMzN3d3d3d3d3d3d3d3d3d3czMzLu7u7u7u7u7u6qqqqqqqqqqqqqqqpmZmaqqqpmZmaqqqpmZmZmZmZmZmXd3d3d3d4iIiHd3d3d3d4iIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiHd3d4iIiHd3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d1VVVWZmZlVVVWZmZlVVVWZmZmZmZnd3d1VVVWZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiHd3d4iIiIiIiIiIiIiIiIiIiHd3d4iIiIiIiIiIiIiIiHd3d4iIiHd3d2ZmZlVVVVVVVVVVVURERERERERERERERDMzM0RERDMzMzMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzM0RERDMzMzMzMzMzM0RERDMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVWZmZlVVVURERGZmZmZmZlVVVWZmZmZmZnd3d3d3d4iIiJmZmXd3d2ZmZnd3d3d3d2ZmZmZmZmZmZnd3d4iIiIiIiIiIiHd3d3d3d4iIiIiIiIiIiIiIiHd3d3d3d5mZmbu7u7u7u5mZmYiIiHd3d6qqqqqqqqqqqpmZmbu7u5mZmWZmZpmZmbu7u5mZmYiIiJmZmbu7u7u7u6qqqru7u7u7u6qqqszMzMzMzMzMzLu7u6qqqpmZmXd3d2ZmZmZmZnd3d3d3d5mZmaqqqpmZmaqqqqqqqpmZmYiIiHd3d3d3d2ZmZpmZmZmZmXd3d2ZmZnd3d4iIiIiIiIiIiHd3d3d3d4iIiIiIiIiIiJmZmYiIiHd3d2ZmZmZmZlVVVWZmZmZmZkRERERERGZmZoiIiHd3d3d3d1VVVURERERERGZmZnd3d3d3d2ZmZnd3d2ZmZmZmZnd3d3d3d3d3d2ZmZlVVVVVVVVVVVWZmZnd3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZnd3d2ZmZlVVVVVVVVVVVWZmZmZmZnd3d3d3d5mZmYiIiHd3d3d3d4iIiGZmZmZmZnd3d3d3d2ZmZlVVVWZmZlVVVVVVVVVVVURERGZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVURERFVVVVVVVURERFVVVURERFVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZlVVVWZmZlVVVVVVVURERERERDMzM0RERERERGZmZmZmZlVVVVVVVXd3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVURERERERERERFVVVURERERERERERERERERERFVVVURERFVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVTMzMzMzMzMzM1VVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d2ZmZlVVVVVVVURERDMzMzMzMzMzM0RERFVVVWZmZlVVVVVVVVVVVWZmZmZmZmZmZnd3d2ZmZmZmZlVVVWZmZlVVVURERERERERERDMzMzMzM0RERFVVVWZmZlVVVVVVVWZmZlVVVURERERERFVVVVVVVVVVVURERERERFVVVVVVVURERERERERERERERERERFVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVURERFVVVURERFVVVVVVVVVVVVVVVWZmZlVVVURERERERERERDMzM1VVVVVVVWZmZmZmZkRERERERERERERERERERERERERERERERERERFVVVTMzM0RERDMzM0RERDMzMyIiIjMzM0RERERERFVVVURERFVVVWZmZlVVVURERERERFVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVURERERERGZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVVVVVWZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d2ZmZnd3d2ZmZmZmZlVVVWZmZmZmZmZmZlVVVVVVVURERFVVVVVVVVVVVWZmZlVVVWZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d1VVVXd3d3d3d2ZmZnd3d4iIiIiIiGZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d2ZmZnd3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d2ZmZnd3d2ZmZmZmZnd3d2ZmZnd3d2ZmZnd3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiHd3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d2ZmZmZmZmZmZnd3d3d3d3d3d2ZmZnd3d3d3d4iIiIiIiJmZmYiIiHd3d4iIiIiIiJmZmYiIiIiIiJmZmYiIiJmZmZmZmYiIiJmZmZmZmZmZmZmZmYiIiHd3d1VVVVVVVURERERERDMzMzMzM0RERERERFVVVURERERERERERERERERERDMzMzMzMzMzMzMzM0RERDMzMzMzM0RERERERERERERERFVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVURERGZmZlVVVVVVVWZmZmZmZlVVVWZmZlVVVWZmZmZmZlVVVVVVVWZmZlVVVWZmZmZmZlVVVVVVVWZmZnd3d2ZmZmZmZlVVVVVVVVVVVURERDMzMzMzMzMzM2ZmZnd3d3d3d1VVVWZmZmZmZpmZmbu7u6qqqoiIiIiIiJmZmYiIiHd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVURERFVVVURERDMzMzMzM0RERGZmZlVVVTMzMzMzM0RERDMzMzMzM0RERDMzM0RERDMzMzMzMzMzM0RERERERERERERERERERERERFVVVVVVVWZmZkRERDMzMzMzM0RERFVVVURERDMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIjMzMzMzM0RERFVVVURERDMzMyIiIiIiIjMzMzMzMzMzMzMzM0RERERERFVVVURERFVVVXd3d2ZmZjMzM0RERHd3d3d3d2ZmZlVVVURERERERERERDMzMzMzMzMzMzMzM0RERDMzMzMzM0RERERERDMzMzMzM0RERGZmZlVVVVVVVWZmZmZmZnd3d3d3d4iIiJmZmaqqqqqqqqqqqpmZmaqqqqqqqqqqqru7u7u7u6qqqpmZmaqqqqqqqpmZmaqqqpmZmXd3d2ZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiHd3d3d3d2ZmZmZmZnd3d2ZmZmZmZlVVVXd3d4iIiHd3d3d3d3d3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERGZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d2ZmZlVVVVVVVWZmZmZmZmZmZmZmZnd3d3d3d2ZmZnd3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiJmZmYiIiHd3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d2ZmZlVVVWZmZnd3d2ZmZnd3d3d3d4iIiIiIiIiIiJmZmZmZmaqqqqqqqszMzN3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7////u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMy7u7u7u7u7u7uqqqqqqqqqqqq7u7uqqqq7u7u7u7vMzMzd3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7d3d3u7u7d3d3d3d3MzMzMzMy7u7u7u7uqqqqqqqqZmZmqqqqZmZmIiIh3d3d3d3d3d3dmZmZVVVVmZmZmZmZ3d3d3d3eIiIiIiIh3d3eIiIiZmZmIiIh3d3eIiIiIiIh3d3d3d3d3d3dmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3eIiIh3d3eIiIh3d3eIiIh3d3d3d3d3d3eIiIiIiIiZmZmZmZmIiIiZmZmZmZmIiIiIiIiIiIh3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVEREREREREREREREQzMzMzMzMzMzMzMzMzMzNERERERERVVVUzMzMzMzNEREREREQzMzNERERVVVVVVVVEREREREREREQzMzMzMzMzMzNEREREREQzMzMzMzNEREQzMzMzMzNEREQzMzMzMzNERERERERVVVVmZmZmZmZERERmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVV3d3d3d3dmZmZ3d3d3d3dmZmZ3d3d3d3d3d3eIiIiIiIhmZmZ3d3eIiIh3d3dmZmZ3d3eZmZmIiIiIiIiZmZnMzMzMzMyqqqqIiIhmZmZ3d3eqqqqqqqqqqqqqqqqIiIhmZma7u7u7u7uZmZmZmZmIiIiZmZm7u7u7u7u7u7u7u7u7u7u7u7vMzMzMzMy7u7u7u7u7u7uIiIh3d3d3d3d3d3eIiIiZmZmqqqqqqqqZmZmZmZl3d3eIiIiIiIhmZmZ3d3eIiIiIiIhmZmZVVVV3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3dmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVV3d3d3d3dmZmZVVVVERERVVVVmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3dVVVVVVVVmZmaIiIhmZmZmZmZmZmZVVVV3d3eIiIhmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVERERERERmZmZ3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3dVVVVVVVVVVVVERERVVVVERERERERVVVVmZmZmZmZmZmZVVVV3d3d3d3d3d3dmZmZmZmZVVVVVVVVERERVVVVVVVVVVVVmZmZVVVVERERVVVVVVVVmZmZmZmZmZmZVVVVmZmZVVVVmZmZVVVVVVVVmZmZVVVVVVVVVVVVEREREREQzMzNERERVVVVVVVVmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVERERERERVVVVERERVVVVERERERERERERERERERERERERERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVEREREREQzMzMzMzNVVVVVVVVmZmZVVVVVVVVmZmZVVVVVVVVVVVVmZmZmZmZ3d3dVVVVVVVVVVVVVVVVEREQzMzNERERVVVVERERVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVEREREREQzMzMzMzMzMzNERERVVVVmZmZVVVVVVVVVVVVVVVVERERVVVVVVVVERERERERVVVVERERVVVVERERVVVVERERERERERERERERVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERVVVV3d3dmZmZVVVVEREREREQzMzNEREREREREREREREREREQzMzNEREQzMzNEREQzMzMzMzNEREQiIiIzMzNVVVVmZmZmZmZVVVV3d3dmZmZVVVVVVVV3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVV3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3eIiIh3d3d3d3d3d3dmZmZmZmZ3d3d3d3dmZmZVVVVmZmZmZmZVVVVmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIiZmZmIiIiZmZmIiIiIiIiIiIiIiIiIiIh3d3eIiIh3d3d3d3d3d3dmZmZ3d3d3d3dmZmZmZmZVVVVmZmZmZmZmZmZ3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZmIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3dmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3eIiIiZmZmIiIiZmZmZmZmIiIiZmZmZmZmZmZmZmZmZmZmZmZmIiIiIiIiIiIh3d3dmZmZVVVVEREQzMzNERERERERVVVVVVVVEREQzMzMzMzNEREQzMzMzMzNEREQzMzMzMzMzMzNERERVVVVVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNERERERERVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVmZmZmZmZmZmZmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVERERVVVVmZmZmZmZVVVVVVVVmZmZVVVVEREQzMzMzMzMiIiIzMzNVVVV3d3eIiIh3d3dmZmZ3d3eIiIi7u7uqqqqqqqqIiIiZmZmZmZmZmZmIiIiIiIhmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVERERERERVVVVmZmZVVVVEREQzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzNERERERERERERVVVVVVVVEREREREQzMzNERERERERmZmZVVVUzMzMzMzMiIiIzMzMiIiIzMzMiIiIiIiIzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzNVVVVEREREREQzMzMiIiIzMzMiIiIiIiIzMzNEREQzMzNERERERERVVVVmZmZ3d3dmZmYzMzNERER3d3d3d3dmZmZVVVVVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzNERERVVVVVVVVVVVVVVVV3d3d3d3eIiIiZmZmZmZmqqqqqqqqqqqqqqqqqqqqqqqqqqqq7u7u7u7uqqqqZmZmqqqq7u7u7u7uqqqqZmZl3d3eIiIh3d3dmZmZ3d3d3d3dmZmZ3d3d3d3d3d3eZmZmZmZl3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3eIiIiIiIh3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3eIiIiIiIiZmZmqqqqqqqqZmZmZmZmZmZmIiIh3d3eIiIh3d3d3d3eIiIh3d3dmZmZ3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3eIiIh3d3dmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3eIiIiZmZmqqqqZmZmqqqq7u7vMzMzd3d3d3d3u7u7////////////////////////////////u7u7///////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////7u7u////7u7u3d3d3d3d3d3d3d3dzMzMu7u7zMzMzMzMzMzMzMzMzMzM3d3dzMzMzMzMzMzMu7u7u7u7u7u7u7u7u7u7u7u7zMzMzMzM3d3dzMzM3d3d3d3d3d3d7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3dzMzMu7u7mZmZmZmZiIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3iIiIiIiIiIiImZmZmZmZiIiIiIiIiIiIiIiIiIiId3d3ZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVZmZmZmZmVVVVZmZmZmZmd3d3d3d3iIiIiIiId3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZmZmZmZmZmZmZmZmZqqqqmZmZqqqqmZmZmZmZiIiId3d3d3d3ZmZmVVVVZmZmVVVVVVVVREREREREREREREREREREREREREREMzMzREREVVVVVVVVVVVVREREREREVVVVREREVVVVVVVVREREREREREREVVVVREREREREVVVVREREREREREREREREREREMzMzREREREREREREREREMzMzVVVVVVVVZmZmVVVVREREREREREREREREZmZmZmZmZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREZmZmZmZmZmZmZmZmZmZmZmZmd3d3iIiIiIiIiIiIiIiId3d3ZmZmZmZmiIiIiIiId3d3d3d3iIiId3d3d3d3mZmZzMzMzMzMqqqqiIiIZmZmZmZmiIiImZmZqqqqiIiIVVVVZmZmu7u7u7u7qqqqqqqqiIiImZmZu7u7zMzMqqqqu7u7u7u7u7u7zMzMu7u7u7u7u7u7u7u7mZmZiIiIiIiIiIiImZmZu7u7qqqqqqqqmZmZiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmZmZmiIiIiIiId3d3iIiId3d3iIiIiIiIiIiIiIiIiIiId3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVREREZmZmZmZmd3d3ZmZmVVVVZmZmVVVVVVVVVVVVZmZmZmZmd3d3ZmZmZmZmZmZmd3d3VVVVVVVVVVVViIiId3d3ZmZmVVVVVVVVZmZmd3d3d3d3ZmZmZmZmZmZmZmZmVVVVREREVVVVVVVVMzMzREREVVVVd3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3ZmZmZmZmZmZmREREVVVVREREREREREREZmZmd3d3ZmZmVVVVZmZmZmZmiIiId3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmVVVVVVVVVVVVZmZmVVVVZmZmVVVVVVVVVVVVREREMzMzREREVVVVZmZmZmZmVVVVVVVVREREZmZmVVVVZmZmVVVVZmZmZmZmVVVVVVVVREREREREREREREREREREREREVVVVREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVZmZmVVVVREREREREREREMzMzMzMzVVVVVVVVVVVVVVVVREREVVVVVVVVZmZmZmZmZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREREREREREREREVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREMzMzREREREREZmZmVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREVVVVREREREREVVVVREREREREREREVVVVZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmREREREREREREREREREREZmZmd3d3ZmZmVVVVREREREREREREREREREREREREREREREREREREMzMzREREMzMzREREMzMzREREMzMzMzMzVVVVZmZmVVVVZmZmd3d3VVVVREREREREVVVVZmZmVVVVVVVVZmZmVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3ZmZmd3d3ZmZmd3d3ZmZmd3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmd3d3d3d3d3d3iIiIZmZmd3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmd3d3d3d3iIiIiIiIiIiIiIiImZmZmZmZmZmZmZmZmZmZmZmZiIiImZmZiIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmd3d3iIiIiIiIiIiIiIiIiIiImZmZmZmZmZmZiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3ZmZmd3d3d3d3ZmZmd3d3ZmZmd3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiImZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZiIiIiIiIiIiId3d3ZmZmZmZmd3d3d3d3d3d3ZmZmVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREZmZmVVVVZmZmZmZmVVVVVVVVREREREREVVVVVVVVVVVVVVVVREREVVVVZmZmZmZmZmZmVVVVVVVVVVVVREREMzMzIiIiMzMzREREVVVVd3d3iIiIiIiIZmZmd3d3d3d3qqqqu7u7u7u7qqqqqqqqqqqqu7u7mZmZiIiId3d3VVVVVVVVZmZmZmZmZmZmd3d3ZmZmZmZmZmZmVVVVVVVVREREREREVVVVVVVVVVVVVVVVMzMzMzMzREREMzMzMzMzREREMzMzMzMzMzMzREREMzMzMzMzMzMzREREMzMzREREREREREREREREMzMzMzMzMzMzMzMzREREZmZmZmZmVVVVMzMzIiIiMzMzMzMzREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzIiIiMzMzREREREREREREREREMzMzIiIiIiIiIiIiIiIiMzMzMzMzMzMzREREREREVVVVZmZmd3d3VVVVMzMzREREd3d3ZmZmZmZmVVVVVVVVZmZmVVVVREREMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVZmZmZmZmd3d3iIiImZmZqqqqmZmZqqqqqqqqu7u7qqqqu7u7qqqqu7u7u7u7u7u7qqqqqqqqqqqqu7u7qqqqqqqqmZmZmZmZiIiIiIiId3d3d3d3ZmZmVVVVd3d3ZmZmZmZmd3d3iIiIiIiIiIiImZmZiIiId3d3d3d3d3d3d3d3d3d3ZmZmiIiIiIiId3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREREREREREREREREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVREREREREZmZmVVVVZmZmd3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVZmZmd3d3d3d3d3d3iIiIiIiImZmZu7u7u7u7u7u7qqqqqqqqqqqqqqqqiIiId3d3d3d3d3d3d3d3iIiIZmZmd3d3ZmZmZmZmZmZmd3d3d3d3d3d3d3d3iIiIiIiId3d3d3d3d3d3d3d3ZmZmd3d3iIiImZmZiIiImZmZqqqqqqqqu7u7u7u7zMzM3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7t3d3d3d3bu7u7u7u7u7u6qqqpmZmaqqqqqqqszMzMzMzMzMzN3d3czMzMzMzMzMzN3d3czMzN3d3czMzN3d3d3d3d3d3d3d3d3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3czMzLu7u6qqqpmZmXd3d2ZmZmZmZnd3d3d3d3d3d4iIiIiIiJmZmZmZmZmZmZmZmYiIiIiIiJmZmYiIiIiIiHd3d3d3d2ZmZmZmZmZmZmZmZlVVVWZmZlVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiHd3d4iIiIiIiIiIiIiIiJmZmYiIiIiIiIiIiIiIiIiIiJmZmYiIiIiIiJmZmZmZmZmZmZmZmZmZmYiIiJmZmYiIiIiIiHd3d3d3d2ZmZlVVVVVVVVVVVVVVVURERFVVVWZmZlVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVWZmZoiIiHd3d2ZmZlVVVURERFVVVVVVVURERDMzM0RERERERERERDMzM0RERERERERERDMzMzMzM0RERERERERERFVVVWZmZmZmZmZmZmZmZnd3d4iIiHd3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVURERFVVVWZmZlVVVXd3d2ZmZmZmZnd3d3d3d3d3d4iIiJmZmXd3d4iIiIiIiIiIiHd3d2ZmZnd3d4iIiKqqqpmZmYiIiHd3d3d3d4iIiLu7u8zMzKqqqpmZmXd3d2ZmZmZmZoiIiJmZmYiIiERERGZmZru7u7u7u6qqqqqqqqqqqoiIiLu7u8zMzLu7u7u7u7u7u6qqqqqqqpmZmaqqqqqqqpmZmYiIiIiIiGZmZnd3d4iIiKqqqru7u6qqqqqqqpmZmZmZmYiIiJmZmXd3d3d3d2ZmZmZmZlVVVWZmZnd3d4iIiIiIiHd3d3d3d3d3d3d3d4iIiIiIiJmZmXd3d3d3d3d3d2ZmZmZmZlVVVVVVVVVVVVVVVURERGZmZmZmZnd3d3d3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVXd3d2ZmZlVVVWZmZlVVVVVVVVVVVVVVVXd3d3d3d1VVVVVVVVVVVWZmZoiIiGZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZkRERERERERERGZmZnd3d3d3d3d3d2ZmZnd3d2ZmZnd3d2ZmZnd3d3d3d3d3d3d3d2ZmZlVVVWZmZlVVVURERERERFVVVXd3d2ZmZlVVVVVVVWZmZnd3d3d3d2ZmZmZmZmZmZlVVVWZmZmZmZlVVVVVVVWZmZlVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZlVVVVVVVVVVVVVVVURERERERFVVVWZmZlVVVVVVVURERERERFVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERERERFVVVURERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERDMzM0RERFVVVVVVVVVVVURERERERFVVVWZmZmZmZmZmZmZmZlVVVWZmZmZmZlVVVVVVVVVVVURERDMzM0RERERERFVVVVVVVURERERERERERFVVVVVVVVVVVVVVVVVVVURERFVVVVVVVURERFVVVURERDMzMzMzMzMzM0RERFVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVURERFVVVURERERERDMzM0RERERERGZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZlVVVURERERERERERFVVVVVVVVVVVVVVVVVVVURERDMzM0RERERERERERERERERERDMzM0RERERERERERERERERERERERDMzMzMzMzMzM0RERDMzM0RERERERFVVVTMzM0RERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d2ZmZnd3d3d3d3d3d3d3d4iIiHd3d4iIiHd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiHd3d4iIiHd3d4iIiHd3d3d3d3d3d2ZmZnd3d3d3d3d3d2ZmZmZmZnd3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d4iIiIiIiIiIiIiIiJmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiIiIiIiIiHd3d4iIiHd3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d4iIiHd3d4iIiIiIiIiIiJmZmZmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiHd3d4iIiIiIiHd3d4iIiIiIiHd3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d3d3d4iIiIiIiIiIiIiIiJmZmZmZmaqqqpmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiJmZmZmZmZmZmYiIiHd3d2ZmZkRERDMzMzMzMzMzMyIiIjMzMzMzM0RERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMzMzM0RERFVVVXd3d2ZmZkRERGZmZnd3d2ZmZlVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVURERERERERERGZmZmZmZmZmZmZmZkRERERERDMzM0RERERERFVVVURERERERERERFVVVWZmZnd3d3d3d2ZmZnd3d6qqqru7u7u7u6qqqqqqqqqqqqqqqoiIiIiIiGZmZlVVVVVVVWZmZmZmZnd3d2ZmZlVVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERERERDMzM0RERDMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMyIiIjMzMzMzM0RERERERDMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM1VVVVVVVURERCIiIiIiIkRERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzM1VVVVVVVWZmZmZmZjMzMyIiIjMzMyIiIjMzMzMzMzMzM0RERERERFVVVXd3d3d3d1VVVTMzM0RERGZmZnd3d2ZmZlVVVVVVVXd3d2ZmZjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERFVVVWZmZnd3d4iIiJmZmaqqqpmZmaqqqqqqqru7u7u7u7u7u6qqqqqqqru7u7u7u5mZmaqqqpmZmaqqqqqqqqqqqpmZmaqqqqqqqoiIiIiIiIiIiIiIiHd3d3d3d2ZmZmZmZmZmZmZmZnd3d3d3d4iIiHd3d3d3d4iIiGZmZnd3d3d3d2ZmZmZmZnd3d3d3d2ZmZmZmZlVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVURERFVVVWZmZlVVVWZmZmZmZmZmZmZmZlVVVURERFVVVURERFVVVVVVVXd3d4iIiKqqqqqqqru7u6qqqszMzLu7u8zMzKqqqpmZmZmZmZmZmXd3d3d3d2ZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZmZmZnd3d4iIiJmZmZmZmZmZmaqqqru7u7u7u7u7u93d3e7u7t3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7d3d27u7u7u7u7u7vMzMy7u7u7u7vMzMzMzMzd3d3d3d3d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMyqqqqZmZmZmZmZmZmqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqZmZmZmZl3d3d3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiZmZmIiIiIiIiIiIiIiIh3d3d3d3eIiIiZmZmIiIh3d3eIiIiIiIiIiIh3d3eIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZVVVVVVVVmZmZ3d3dmZmZVVVVEREREREQzMzMzMzNEREQzMzNERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZVVVV3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3dmZmZmZmZmZmZERERVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVmZmZ3d3d3d3eIiIh3d3dmZmZ3d3d3d3d3d3d3d3eZmZmIiIh3d3eIiIiIiIh3d3d3d3dmZmaZmZm7u7uqqqqIiIiZmZmIiIiIiIi7u7vMzMyqqqqZmZmIiIh3d3dmZmZ3d3d3d3dmZmZERERmZma7u7vMzMy7u7u7u7uqqqqqqqqqqqq7u7u7u7uqqqqZmZmZmZmIiIiZmZmIiIiZmZmIiIiIiIh3d3d3d3d3d3eIiIiZmZmZmZmqqqqZmZmZmZl3d3eIiIiIiIh3d3dmZmZ3d3d3d3dVVVVVVVV3d3d3d3d3d3d3d3d3d3dVVVV3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVmZmZ3d3d3d3dmZmZERERERERVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVERERVVVVmZmZmZmZVVVVVVVVERERVVVV3d3d3d3eIiIhmZmZVVVVVVVVVVVVmZmZVVVVVVVVERERERERERERmZmZ3d3d3d3d3d3dmZmZ3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZ3d3d3d3dVVVVERERERERmZmZ3d3dmZmZVVVVERERVVVVmZmZmZmZVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVEREQzMzNVVVVmZmZmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZERERVVVVERERVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVERERERERERERERERERERVVVVERERERERVVVVVVVVERERVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVEREREREREREQzMzMiIiJERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3eIiIhmZmZVVVVEREQzMzNERERERERVVVVmZmZmZmZVVVVVVVVEREREREREREREREREREREREREREREREREREREREREREREREREREQzMzMiIiIzMzMzMzNEREREREREREQzMzNEREQzMzNERERERERERERERERVVVVERERERERVVVVERERVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVERERERERERERERERERERERERVVVVERERVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZVVVVmZmZmZmZmZmZmZmZ3d3d3d3dmZmZ3d3d3d3eIiIh3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIiZmZmIiIh3d3eIiIh3d3eIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZmZmZmZmZVVVVmZmZmZmZmZmZ3d3d3d3d3d3d3d3eIiIiIiIiIiIiZmZmIiIiZmZmIiIiZmZmIiIiZmZmIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3eIiIh3d3d3d3d3d3dmZmZ3d3dmZmZmZmZ3d3d3d3d3d3eIiIh3d3eIiIiIiIiIiIiZmZmIiIiIiIiIiIiIiIiIiIiIiIiZmZmIiIiIiIiZmZmIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIiZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmIiIh3d3dVVVUzMzMzMzMiIiIiIiIiIiIzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzNERERVVVVmZmZVVVVERERVVVV3d3dmZmZmZmZVVVVVVVVVVVVVVVVmZmZVVVVERERERERERERVVVVERERERERERERVVVVVVVV3d3dmZmZVVVVEREQzMzMzMzMzMzNERERVVVVERERERERERERERERERERVVVV3d3dmZmZmZmZVVVWIiIi7u7u7u7uqqqqqqqqqqqqqqqqqqqqZmZl3d3dmZmZmZmZmZmZ3d3d3d3dmZmZVVVVERERVVVVVVVVmZmZVVVVEREQzMzMzMzNERERVVVVEREQzMzMzMzMzMzMzMzNEREREREQzMzNEREQzMzMzMzMzMzMiIiJEREREREQzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzNEREQzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMiIiIzMzNERERVVVVVVVVVVVVVVVUzMzMzMzMiIiIzMzMzMzMzMzMzMzNERERVVVVmZmaZmZmZmZlmZmYzMzNERER3d3d3d3dVVVVVVVVERERmZmZVVVVEREQzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERVVVVmZmaIiIiIiIiZmZmZmZmqqqqqqqqZmZmqqqqqqqq7u7uqqqqqqqqqqqqqqqqqqqqqqqqZmZmqqqqqqqqqqqqZmZmZmZmZmZmIiIiIiIiIiIiZmZmZmZmIiIiIiIh3d3dmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVmZmZVVVVmZmZVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVERERERERERERVVVVVVVVVVVVmZmZ3d3eIiIiqqqq7u7u7u7vMzMy7u7u7u7uqqqqqqqqZmZmIiIh3d3dmZmZmZmZmZmZ3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3dVVVVmZmZmZmZ3d3eZmZmIiIiZmZmZmZm7u7u7u7vMzMzMzMzd3d3d3d3d3d3u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d7u7u3d3d7u7u3d3d3d3d3d3d7u7u3d3d3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzMzMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMu7u7u7u7zMzMqqqqmZmZd3d3iIiIiIiId3d3d3d3d3d3VVVVZmZmVVVVVVVVZmZmZmZmZmZmd3d3d3d3iIiIiIiId3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZiIiIiIiId3d3iIiId3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVREREVVVVREREVVVVVVVVREREZmZmZmZmVVVVZmZmd3d3ZmZmZmZmZmZmd3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVREREREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3mZmZiIiId3d3d3d3d3d3ZmZmd3d3ZmZmZmZmVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVZmZmZmZmiIiImZmZiIiId3d3d3d3ZmZmZmZmd3d3mZmZd3d3d3d3d3d3iIiId3d3d3d3ZmZmd3d3qqqqqqqqmZmZmZmZiIiIiIiIqqqqu7u7u7u7qqqqmZmZZmZmVVVVd3d3d3d3VVVVZmZmd3d3zMzMu7u7u7u7qqqqu7u7qqqqmZmZmZmZqqqqmZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3ZmZmZmZmd3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmd3d3ZmZmiIiId3d3d3d3ZmZmd3d3d3d3d3d3d3d3ZmZmZmZmd3d3d3d3d3d3ZmZmVVVVVVVVVVVVZmZmZmZmd3d3iIiIVVVVVVVVVVVVREREREREVVVVZmZmZmZmZmZmZmZmZmZmREREREREVVVVREREVVVVZmZmVVVVREREREREVVVVVVVVZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVREREREREREREZmZmd3d3iIiIZmZmd3d3iIiIiIiIiIiId3d3d3d3ZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVREREZmZmd3d3ZmZmVVVVZmZmVVVVZmZmZmZmZmZmZmZmd3d3d3d3VVVVVVVVVVVVVVVVVVVVREREREREVVVVZmZmd3d3d3d3ZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVREREREREMzMzREREVVVVZmZmZmZmVVVVREREVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREREREREREREREREREREREREREREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREVVVVVVVVZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3ZmZmVVVVZmZmVVVVVVVVREREREREMzMzREREREREVVVVVVVVVVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREMzMzMzMzREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVREREREREREREREREREREZmZmZmZmZmZmZmZmVVVVZmZmVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3VVVVVVVVREREREREREREVVVVZmZmZmZmVVVVVVVVREREREREREREREREREREVVVVREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzREREREREVVVVREREREREREREMzMzREREREREVVVVVVVVREREMzMzREREMzMzREREREREREREREREREREMzMzMzMzREREVVVVREREREREMzMzREREREREREREZmZmZmZmREREREREREREREREREREREREREREREREVVVVZmZmVVVVVVVVZmZmZmZmd3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmd3d3ZmZmd3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiImZmZiIiIiIiIiIiImZmZiIiIiIiId3d3iIiId3d3d3d3d3d3ZmZmZmZmd3d3d3d3ZmZmZmZmVVVVZmZmZmZmZmZmZmZmd3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiImZmZiIiImZmZmZmZmZmZiIiImZmZiIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3ZmZmZmZmd3d3d3d3ZmZmZmZmZmZmd3d3d3d3d3d3d3d3iIiIiIiIiIiImZmZiIiImZmZmZmZmZmZqqqqmZmZmZmZmZmZiIiIiIiIiIiIiIiIiIiIiIiId3d3iIiId3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZiIiImZmZmZmZmZmZmZmZqqqqmZmZmZmZmZmZmZmZmZmZmZmZiIiId3d3ZmZmREREREREMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzIiIiMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzZmZmVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREVVVVREREREREREREREREd3d3iIiIZmZmVVVVMzMzMzMzIiIiMzMzMzMzREREREREREREREREREREREREREREVVVVZmZmZmZmVVVVREREZmZmmZmZu7u7qqqqmZmZqqqqqqqqqqqqqqqqiIiIZmZmVVVVZmZmd3d3d3d3ZmZmREREVVVVVVVVZmZmVVVVZmZmVVVVREREMzMzREREZmZmREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREVVVVVVVVREREMzMzMzMzREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzVVVVZmZmVVVVREREREREREREMzMzMzMzREREMzMzREREZmZmiIiIiIiImZmZiIiIZmZmREREMzMzd3d3d3d3VVVVVVVVVVVVREREREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzREREMzMzMzMzMzMzREREVVVVVVVVVVVViIiIiIiImZmZqqqqqqqqmZmZiIiImZmZqqqqqqqqu7u7qqqqqqqqqqqqmZmZqqqqqqqqqqqqqqqqqqqqmZmZmZmZmZmZmZmZmZmZiIiIiIiImZmZiIiId3d3ZmZmZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVZmZmVVVVREREREREREREVVVVZmZmZmZmZmZmiIiIqqqqu7u7zMzMu7u7zMzMqqqqqqqqqqqqmZmZiIiIZmZmZmZmd3d3iIiId3d3d3d3ZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmd3d3d3d3ZmZmZmZmZmZmd3d3iIiImZmZqqqqqqqqqqqqu7u7zMzMzMzM3d3d3d3d7u7u////7u7u////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3e7u7u7u7t3d3d3d3d3d3czMzN3d3czMzKqqqpmZmZmZmYiIiIiIiGZmZlVVVVVVVVVVVVVVVWZmZnd3d2ZmZnd3d3d3d3d3d4iIiIiIiIiIiJmZmYiIiIiIiJmZmYiIiHd3d4iIiIiIiIiIiIiIiHd3d4iIiIiIiIiIiIiIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiHd3d2ZmZmZmZmZmZlVVVVVVVVVVVURERERERERERERERERERDMzMzMzMzMzM0RERERERERERFVVVVVVVWZmZnd3d2ZmZlVVVURERERERFVVVVVVVVVVVURERERERERERERERDMzM0RERERERERERERERERERERERFVVVVVVVWZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d2ZmZoiIiIiIiHd3d3d3d4iIiIiIiHd3d4iIiIiIiHd3d3d3d2ZmZmZmZmZmZmZmZnd3d2ZmZmZmZlVVVURERFVVVWZmZmZmZmZmZmZmZlVVVWZmZnd3d3d3d4iIiJmZmYiIiHd3d2ZmZlVVVWZmZoiIiHd3d3d3d4iIiJmZmZmZmYiIiHd3d3d3d4iIiJmZmaqqqpmZmYiIiHd3d5mZmbu7u6qqqqqqqoiIiFVVVVVVVYiIiHd3d1VVVVVVVXd3d7u7u8zMzKqqqqqqqqqqqqqqqnd3d2ZmZoiIiJmZmYiIiIiIiJmZmXd3d3d3d4iIiHd3d2ZmZmZmZmZmZmZmZoiIiIiIiIiIiHd3d4iIiIiIiHd3d3d3d3d3d3d3d3d3d4iIiGZmZmZmZnd3d3d3d3d3d4iIiIiIiHd3d1VVVVVVVVVVVWZmZmZmZnd3d2ZmZmZmZlVVVVVVVWZmZlVVVVVVVURERERERFVVVWZmZnd3d1VVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVURERERERDMzMzMzM0RERGZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVURERFVVVURERERERERERGZmZnd3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZlVVVURERFVVVURERERERERERFVVVWZmZmZmZnd3d2ZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZlVVVVVVVURERERERFVVVVVVVURERERERGZmZnd3d2ZmZmZmZmZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZlVVVURERERERDMzM0RERERERFVVVWZmZmZmZmZmZlVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZlVVVWZmZlVVVVVVVURERERERDMzM0RERDMzM0RERDMzM0RERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVWZmZmZmZlVVVWZmZmZmZmZmZnd3d3d3d3d3d3d3d2ZmZnd3d2ZmZmZmZlVVVURERFVVVURERDMzM1VVVVVVVVVVVVVVVURERFVVVVVVVURERFVVVURERFVVVURERERERFVVVURERFVVVURERERERDMzMzMzM0RERFVVVXd3d1VVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZlVVVWZmZlVVVWZmZlVVVURERDMzM1VVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZkRERERERERERGZmZmZmZmZmZmZmZkRERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVTMzMzMzMzMzM0RERERERFVVVWZmZlVVVVVVVWZmZlVVVURERERERERERERERERERERERDMzMzMzM0RERDMzM0RERERERERERERERERERERERFVVVURERERERERERGZmZlVVVVVVVXd3d2ZmZlVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZnd3d3d3d4iIiHd3d3d3d3d3d3d3d3d3d4iIiHd3d5mZmZmZmZmZmYiIiJmZmZmZmYiIiJmZmYiIiIiIiIiIiJmZmYiIiHd3d4iIiGZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d4iIiHd3d4iIiJmZmYiIiJmZmYiIiJmZmYiIiJmZmZmZmYiIiIiIiHd3d4iIiHd3d4iIiHd3d4iIiHd3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiIiIiJmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiIiIiIiIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiHd3d4iIiIiIiJmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiJmZmYiIiIiIiIiIiGZmZmZmZlVVVVVVVURERERERDMzMzMzMyIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERDMzM1VVVYiIiGZmZlVVVURERFVVVWZmZlVVVURERERERERERFVVVURERFVVVURERERERDMzM0RERERERDMzMyIiIlVVVYiIiHd3d0RERDMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERDMzMzMzM0RERERERFVVVVVVVVVVVURERGZmZqqqqru7u6qqqqqqqpmZmaqqqqqqqqqqqoiIiHd3d2ZmZnd3d2ZmZlVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVTMzM0RERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM0RERDMzM0RERFVVVVVVVURERERERDMzM0RERERERERERDMzM0RERDMzMzMzMzMzMzMzM0RERFVVVVVVVVVVVVVVVURERERERERERERERDMzM0RERIiIiLu7u4iIiGZmZnd3d2ZmZjMzMzMzM2ZmZmZmZmZmZlVVVURERERERERERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVWZmZnd3d3d3d4iIiIiIiJmZmYiIiIiIiHd3d4iIiIiIiJmZmaqqqqqqqru7u6qqqqqqqqqqqqqqqqqqqqqqqoiIiJmZmYiIiJmZmZmZmYiIiIiIiIiIiJmZmYiIiHd3d2ZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVWZmZmZmZlVVVWZmZmZmZmZmZmZmZlVVVURERERERERERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d6qqqru7u7u7u7u7u6qqqqqqqqqqqqqqqpmZmXd3d2ZmZmZmZnd3d3d3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVXd3d3d3d4iIiHd3d3d3d3d3d4iIiJmZmaqqqqqqqru7u7u7u8zMzN3d3d3d3d3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3u7u7d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3MzMy7u7u7u7uZmZl3d3dmZmZmZmZmZmZmZmZVVVVVVVVmZmZ3d3d3d3d3d3eIiIiZmZmIiIiZmZmZmZmZmZmZmZmIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiZmZmIiIiIiIiZmZmIiIh3d3d3d3d3d3dmZmZVVVVERERERERERERVVVVVVVVEREREREREREQzMzNEREQzMzMzMzMiIiIzMzMzMzMzMzNERERERERERERERERERERVVVVEREREREREREQzMzNEREQzMzNEREREREQzMzMzMzNERERERERERERERERERERmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3eIiIiIiIh3d3d3d3dmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVmZmZmZmZmZmZVVVVVVVVERERERERVVVV3d3d3d3dmZmZmZmZVVVV3d3eIiIiIiIiZmZmZmZmZmZl3d3dmZmZ3d3dmZmZ3d3d3d3d3d3eZmZm7u7uqqqqIiIh3d3eZmZmZmZmZmZmZmZmZmZmIiIiIiIiZmZmqqqqqqqqIiIh3d3dVVVVmZmZ3d3d3d3dVVVVVVVVmZmaqqqq7u7uqqqqIiIiZmZmqqqqIiIh3d3d3d3eZmZmqqqqqqqqIiIh3d3d3d3eIiIh3d3d3d3dmZmZ3d3dmZmZ3d3eZmZmIiIh3d3d3d3d3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZ3d3eIiIh3d3dmZmZVVVVVVVVERERVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVmZmZmZmZVVVVERERmZmZVVVVVVVVVVVVVVVVERERVVVVVVVVEREREREREREQzMzNERERVVVVVVVVmZmZmZmZVVVVERERmZmZmZmZ3d3dmZmZ3d3dmZmZVVVVVVVVVVVVVVVVVVVVERERVVVVmZmZ3d3dmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVERERERERERERVVVVVVVVmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERERERVVVVmZmZ3d3dmZmZmZmZ3d3dmZmZ3d3d3d3dmZmZ3d3dmZmZmZmZVVVVVVVVERERERERERERERERVVVV3d3dmZmZVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVERERERERERERERERERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERmZmZmZmZmZmZVVVVmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZVVVVERERERERERERERERmZmZVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERmZmZ3d3dmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVERERERERVVVVVVVVmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZVVVVmZmZmZmZmZmZ3d3d3d3eIiIh3d3d3d3dVVVVVVVVERERVVVVVVVVmZmZ3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVEREQzMzMzMzNERERVVVVERERVVVVERERVVVVVVVVVVVVVVVVEREREREREREREREREREQzMzMzMzMzMzMzMzNERERERERVVVVVVVVVVVVERERVVVVVVVVERERVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVV3d3d3d3dmZmZ3d3dmZmZmZmZmZmZmZmZ3d3d3d3eIiIh3d3d3d3dmZmZ3d3d3d3dmZmZ3d3eIiIh3d3d3d3d3d3eIiIiIiIiIiIiZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmIiIiIiIh3d3d3d3d3d3dmZmZmZmZmZmZVVVVmZmZmZmZVVVVmZmZmZmZmZmZ3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIiZmZmZmZmZmZmIiIiZmZmIiIiZmZmIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3dmZmZmZmZmZmZ3d3dmZmZ3d3dmZmaIiIh3d3eIiIiIiIiIiIiIiIiIiIiZmZmIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZmIiIiIiIh3d3eIiIh3d3eIiIh3d3eIiIiZmZmIiIiIiIiIiIiIiIiZmZmIiIiIiIiIiIiZmZmZmZmIiIiIiIh3d3dmZmZ3d3dVVVVVVVVEREREREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNERERmZmZVVVVVVVVERERVVVVVVVVERERERERERERVVVVERERVVVVVVVVEREQzMzMiIiIzMzMzMzMiIiIzMzNVVVVmZmZVVVVVVVVEREREREREREQzMzNERERERERERERVVVVEREREREREREQzMzMzMzMzMzMzMzNERERVVVVVVVVERERERER3d3e7u7u7u7uqqqqqqqqZmZmqqqqqqqqZmZmIiIhmZmZ3d3dmZmZVVVVVVVVmZmZVVVVVVVVVVVVmZmZmZmZEREQzMzNEREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzMzMzMiIiIzMzMzMzMzMzNEREQzMzNERERERERERERERERERERERERERERVVVVVVVVVVVVEREREREREREREREQzMzNEREQzMzNERERERERERERERERERERmZmZmZmZVVVVVVVVVVVVERERERERERERERERVVVV3d3eZmZlmZmZERERVVVV3d3dVVVUzMzNmZmZmZmZVVVVVVVVVVVVEREREREREREQzMzNEREQzMzMzMzMzMzMzMzMiIiIiIiIzMzNERERVVVVmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmaIiIiIiIiZmZmqqqqqqqqZmZmqqqqqqqqqqqqqqqqZmZmZmZmZmZmZmZmZmZmIiIiZmZmIiIiIiIiIiIiIiIiIiIh3d3dmZmZmZmZmZmZmZmZVVVVVVVVmZmZ3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZERERVVVVERERVVVVVVVVVVVVmZmZVVVVERERVVVVVVVVERERVVVVERERVVVVVVVVERERERERERERVVVVVVVV3d3d3d3d3d3d3d3dVVVVERERVVVVERERERERVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmaIiIiZmZmqqqqqqqqqqqqqqqqqqqqqqqqIiIh3d3d3d3d3d3d3d3d3d3dVVVVERERVVVVVVVVmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3eIiIiIiIiZmZmZmZmqqqq7u7u7u7vMzMzMzMzMzMzd3d3MzMzd3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzM3d3d3d3d7u7u3d3d7u7u3d3d7u7u7u7u3d3d7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMu7u7qqqqmZmZiIiIiIiIiIiIiIiIiIiIiIiImZmZmZmZiIiImZmZmZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3iIiIiIiIiIiImZmZmZmZmZmZiIiImZmZiIiId3d3ZmZmZmZmZmZmZmZmREREREREMzMzMzMzMzMzIiIiMzMzVVVVMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzREREMzMzREREMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3iIiIiIiIiIiId3d3d3d3ZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREVVVVZmZmiIiIZmZmVVVVVVVVVVVViIiImZmZmZmZmZmZqqqqiIiIZmZmZmZmiIiId3d3d3d3d3d3iIiImZmZmZmZmZmZiIiImZmZqqqqqqqqqqqqiIiImZmZmZmZiIiIiIiImZmZmZmZiIiId3d3VVVVZmZmd3d3ZmZmVVVVZmZmd3d3iIiIqqqqmZmZiIiIiIiIiIiIiIiId3d3ZmZmmZmZqqqqmZmZd3d3d3d3d3d3d3d3d3d3iIiId3d3ZmZmZmZmd3d3mZmZiIiId3d3d3d3ZmZmd3d3d3d3d3d3d3d3VVVVZmZmd3d3ZmZmZmZmZmZmVVVVd3d3d3d3d3d3ZmZmVVVVVVVVREREVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVZmZmZmZmZmZmVVVVVVVVZmZmVVVVVVVVVVVVREREVVVVVVVVREREVVVVREREMzMzREREVVVVZmZmZmZmVVVVVVVVZmZmZmZmZmZmZmZmd3d3ZmZmZmZmd3d3ZmZmZmZmVVVVZmZmZmZmVVVVZmZmd3d3d3d3d3d3ZmZmZmZmZmZmd3d3d3d3ZmZmZmZmd3d3ZmZmVVVVVVVVVVVVREREREREREREVVVVZmZmd3d3d3d3ZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmd3d3ZmZmZmZmd3d3ZmZmZmZmd3d3ZmZmZmZmd3d3ZmZmZmZmVVVVVVVVREREREREREREVVVVd3d3ZmZmZmZmVVVVZmZmd3d3ZmZmd3d3ZmZmd3d3d3d3d3d3d3d3ZmZmZmZmVVVVREREVVVVREREVVVVREREREREREREREREVVVVVVVVREREVVVVVVVVVVVVZmZmZmZmVVVVVVVVREREREREREREVVVVZmZmd3d3ZmZmVVVVZmZmZmZmd3d3d3d3ZmZmZmZmd3d3d3d3d3d3d3d3ZmZmZmZmVVVVREREREREVVVVVVVVVVVVVVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVREREMzMzREREREREZmZmd3d3ZmZmVVVVVVVVZmZmZmZmZmZmVVVVZmZmVVVVd3d3ZmZmZmZmZmZmZmZmVVVVVVVVREREREREZmZmd3d3d3d3ZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3ZmZmREREREREREREVVVVd3d3d3d3ZmZmZmZmd3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREMzMzMzMzREREVVVVVVVVVVVVREREREREREREREREREREREREVVVVVVVVREREREREMzMzREREMzMzREREREREMzMzREREREREVVVVREREZmZmVVVVZmZmd3d3iIiId3d3d3d3VVVVREREVVVVVVVVREREVVVVVVVVREREVVVVZmZmVVVVVVVVVVVVZmZmVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiIiIiImZmZmZmZmZmZqqqqmZmZmZmZiIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmd3d3d3d3ZmZmZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmd3d3d3d3d3d3iIiIiIiIiIiImZmZiIiImZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZiIiIiIiId3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiIZmZmd3d3ZmZmd3d3iIiId3d3d3d3iIiIiIiIiIiIiIiIiIiImZmZmZmZiIiImZmZmZmZmZmZmZmZiIiIiIiIiIiIiIiIiIiId3d3iIiId3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZiIiIiIiIiIiImZmZiIiIiIiId3d3d3d3ZmZmZmZmZmZmVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzVVVVREREREREREREVVVVREREMzMzREREREREMzMzREREMzMzIiIiERERERERIiIiMzMzMzMzREREVVVVVVVVREREVVVVZmZmZmZmVVVVMzMzMzMzMzMzREREREREREREREREREREIiIiIiIiIiIiMzMzREREREREREREREREREREVVVVmZmZu7u7u7u7qqqqqqqqqqqqmZmZqqqqmZmZd3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmREREREREREREVVVVVVVVREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzREREMzMzREREMzMzREREREREMzMzREREVVVVVVVVREREMzMzMzMzREREREREREREREREREREREREREREREREVVVVZmZmZmZmVVVVVVVVVVVVREREREREREREREREVVVViIiIiIiIVVVVVVVVZmZmd3d3VVVVMzMzZmZmd3d3ZmZmVVVVVVVVREREREREREREREREREREMzMzVVVVREREMzMzMzMzREREREREVVVVVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3iIiImZmZmZmZiIiIiIiIiIiImZmZmZmZmZmZmZmZmZmZmZmZmZmZiIiIiIiIiIiImZmZmZmZiIiIiIiIZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVVVVVREREREREVVVVVVVVVVVVREREVVVVVVVVREREVVVVVVVVREREVVVVREREVVVVREREVVVVREREREREVVVVVVVVVVVVREREREREVVVVREREREREREREVVVVVVVVd3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVZmZmZmZmZmZmiIiImZmZmZmZqqqqqqqqmZmZiIiIiIiIiIiIiIiIZmZmZmZmVVVVVVVVVVVVZmZmd3d3d3d3d3d3d3d3d3d3iIiImZmZiIiImZmZmZmZqqqqqqqqu7u7u7u7zMzMzMzMzMzMzMzMzMzMzMzM7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7t3d3d3d3czMzN3d3d3d3d3d3e7u7u7u7t3d3e7u7t3d3d3d3e7u7t3d3e7u7t3d3d3d3e7u7t3d3d3d3d3d3czMzN3d3bu7u8zMzLu7u7u7u8zMzMzMzMzMzMzMzN3d3czMzMzMzMzMzMzMzLu7u7u7u7u7u6qqqqqqqpmZmZmZmYiIiJmZmYiIiIiIiIiIiHd3d3d3d3d3d4iIiIiIiIiIiJmZmYiIiIiIiHd3d4iIiIiIiHd3d4iIiIiIiHd3d2ZmZlVVVVVVVURERERERERERERERERERERERERERDMzM0RERDMzMyIiIjMzMyIiIjMzMzMzMzMzMyIiIjMzMyIiIiIiIjMzMyIiIiIiIjMzM0RERERERERERERERERERERERERERERERERERERERERERERERFVVVWZmZlVVVWZmZmZmZmZmZnd3d3d3d2ZmZnd3d3d3d2ZmZmZmZmZmZmZmZnd3d2ZmZmZmZnd3d3d3d4iIiIiIiIiIiIiIiIiIiHd3dwD//wAAiIiId3d3ZmZmZmZmZmZmVVVVZmZmVVVVVVVVREREREREREREREREVVVVVVVVREREVVVVVVVVVVVVREREREREVVVVZmZmVVVVZmZmd3d3ZmZmZmZmZmZmZmZmiIiImZmZiIiIiIiImZmZiIiId3d3d3d3iIiId3d3iIiImZmZmZmZmZmZiIiId3d3iIiIqqqqu7u7zMzMqqqqmZmZmZmZqqqqd3d3d3d3iIiIiIiIiIiIZmZmZmZmZmZmiIiIiIiIZmZmd3d3ZmZmd3d3qqqqmZmZiIiImZmZiIiId3d3ZmZmVVVVd3d3iIiIiIiId3d3ZmZmZmZmZmZmd3d3iIiIZmZmZmZmZmZmZmZmd3d3mZmZd3d3ZmZmVVVVVVVVZmZmd3d3ZmZmVVVVZmZmZmZmZmZmd3d3iIiIZmZmd3d3d3d3ZmZmVVVVREREREREVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmiIiIiIiId3d3ZmZmd3d3ZmZmZmZmZmZmZmZmVVVVREREREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmREREVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmd3d3iIiId3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3ZmZmVVVVZmZmVVVVZmZmZmZmd3d3ZmZmd3d3ZmZmVVVVVVVVZmZmZmZmVVVVVVVVZmZmd3d3d3d3d3d3ZmZmZmZmZmZmd3d3ZmZmd3d3d3d3d3d3ZmZmZmZmZmZmVVVVVVVVREREZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmVVVVREREREREREREREREVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmZmZmd3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3ZmZmZmZmVVVVZmZmVVVVVVVVZmZmZmZmVVVVREREREREVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVZmZmd3d3ZmZmVVVVVVVVZmZmVVVVZmZmZmZmVVVVZmZmZmZmd3d3ZmZmZmZmZmZmZmZmREREVVVVZmZmd3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3iIiId3d3ZmZmREREVVVVVVVVd3d3iIiId3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVREREVVVVREREMzMzMzMzREREVVVVVVVVZmZmVVVVVVVVREREREREVVVVVVVVVVVVVVVVREREREREREREREREREREREREREREMzMzREREREREMzMzREREREREVVVVVVVVVVVVZmZmZmZmd3d3VVVVVVVVREREVVVVREREREREREREVVVVREREVVVVVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmVVVVVVVVZmZmVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVZmZmVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmd3d3d3d3mZmZiIiImZmZiIiIiIiId3d3d3d3d3d3d3d3ZmZmd3d3iIiId3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3iIiIiIiImZmZmZmZmZmZmZmZmZmZmZmZmZmZiIiImZmZiIiImZmZiIiIiIiId3d3iIiId3d3d3d3d3d3d3d3ZmZmZmZmZmZmVVVVZmZmZmZmd3d3d3d3d3d3iIiIiIiImZmZiIiIiIiIiIiImZmZiIiImZmZmZmZmZmZiIiIiIiIiIiIiIiIiIiId3d3d3d3iIiImZmZiIiId3d3ZmZmd3d3d3d3d3d3iIiIZmZmZmZmd3d3ZmZmd3d3d3d3iIiIiIiImZmZmZmZmZmZqqqqqqqqmZmZmZmZmZmZmZmZiIiIiIiId3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3iIiId3d3d3d3d3d3d3d3d3d3ZmZmZmZmVVVVVVVVREREREREREREREREREREREREVVVVREREMzMzREREREREREREREREMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiREREMzMzREREREREREREREREVVVVZmZmd3d3d3d3ZmZmREREREREREREREREVVVVREREREREMzMzMzMzMzMzMzMzREREREREREREVVVVREREMzMzVVVVqqqqu7u7u7u7qqqqmZmZmZmZmZmZmZmZiIiId3d3ZmZmVVVVVVVVVVVVZmZmZmZmVVVVVVVVZmZmd3d3VVVVMzMzVVVVREREREREREREREREMzMzREREREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzREREMzMzREREMzMzREREREREREREREREREREREREREREREREREREREREMzMzMzMzREREMzMzREREREREREREVVVVVVVVVVVVZmZmd3d3d3d3ZmZmZmZmVVVVREREVVVVVVVVREREZmZmZmZmZmZmVVVVZmZmd3d3d3d3REREREREd3d3d3d3ZmZmZmZmZmZmVVVVREREREREREREREREMzMzREREREREREREMzMzREREVVVVZmZmVVVVZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmd3d3iIiIiIiIiIiId3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3iIiImZmZiIiId3d3ZmZmREREVVVVVVVVVVVVVVVVVVVVREREVVVVZmZmVVVVREREVVVVREREREREREREREREREREVVVVVVVVVVVVREREREREREREREREVVVVREREREREVVVVVVVVREREREREVVVVREREVVVVREREVVVVREREREREREREREREREREREREREREVVVVZmZmVVVVZmZmZmZmVVVVZmZmd3d3ZmZmZmZmd3d3d3d3d3d3d3d3ZmZmZmZmVVVVZmZmZmZmZmZmiIiImZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZd3d3ZmZmVVVVVVVVZmZmd3d3d3d3d3d3d3d3d3d3iIiIiIiImZmZmZmZqqqqu7u7u7u7u7u7u7u7zMzMzMzMu7u7qqqqu7u7zMzM7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////+7u7v///+7u7u7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3e7u7t3d3d3d3d3d3d3d3czMzLu7u7u7u7u7u7u7u6qqqru7u7u7u7u7u8zMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzKqqqqqqqpmZmYiIiHd3d3d3d3d3d3d3d4iIiIiIiIiIiJmZmaqqqqqqqpmZmZmZmYiIiHd3d2ZmZmZmZlVVVVVVVURERERERERERERERCIiIjMzMzMzMzMzMyIiIjMzMzMzM0RERDMzM0RERERERFVVVURERERERERERDMzMzMzM0RERERERERERDMzMzMzM0RERDMzMzMzM0RERFVVVVVVVVVVVWZmZlVVVVVVVWZmZlVVVVVVVWZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZoiIiHd3d4iIiIiIiIiIiIiIiIiIiHd3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVURERGZmZlVVVVVVVVVVVVVVVVVVVURERFVVVXd3d2ZmZlVVVVVVVWZmZmZmZmZmZmZmZnd3d2ZmZmZmZnd3d4iIiJmZmYiIiIiIiHd3d4iIiIiIiHd3d4iIiIiIiIiIiJmZmZmZmZmZmaqqqoiIiIiIiKqqqszMzMzMzKqqqqqqqqqqqoiIiGZmZlVVVVVVVWZmZnd3d2ZmZmZmZmZmZqqqqru7u4iIiHd3d2ZmZmZmZoiIiJmZmaqqqoiIiIiIiGZmZlVVVVVVVWZmZnd3d4iIiHd3d2ZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZnd3d3d3d4iIiGZmZlVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZnd3d5mZmYiIiHd3d2ZmZmZmZmZmZkRERERERERERFVVVVVVVVVVVVVVVURERFVVVWZmZnd3d5mZmYiIiGZmZmZmZmZmZmZmZnd3d2ZmZmZmZkRERERERERERERERGZmZmZmZoiIiHd3d3d3d2ZmZlVVVVVVVURERERERGZmZlVVVURERERERFVVVWZmZnd3d2ZmZnd3d3d3d2ZmZoiIiJmZmYiIiIiIiGZmZmZmZnd3d3d3d2ZmZmZmZmZmZmZmZnd3d3d3d3d3d2ZmZnd3d3d3d3d3d2ZmZmZmZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d4iIiHd3d3d3d3d3d2ZmZnd3d2ZmZnd3d2ZmZnd3d2ZmZnd3d3d3d3d3d3d3d2ZmZmZmZnd3d4iIiIiIiHd3d2ZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZnd3d3d3d3d3d3d3d3d3d2ZmZlVVVWZmZlVVVTMzM0RERERERERERFVVVVVVVVVVVVVVVXd3d2ZmZmZmZlVVVVVVVVVVVXd3d3d3d3d3d2ZmZlVVVVVVVVVVVWZmZnd3d2ZmZmZmZmZmZmZmZnd3d3d3d3d3d2ZmZlVVVWZmZnd3d4iIiHd3d1VVVVVVVURERERERERERERERFVVVURERFVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVURERFVVVXd3d4iIiHd3d2ZmZlVVVVVVVURERFVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVXd3d3d3d4iIiIiIiHd3d3d3d3d3d1VVVWZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZnd3d4iIiIiIiIiIiIiIiHd3d1VVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERDMzM0RERFVVVWZmZmZmZlVVVURERERERFVVVVVVVWZmZlVVVURERERERFVVVURERERERERERDMzM0RERERERERERDMzM0RERERERERERFVVVVVVVVVVVURERFVVVURERFVVVURERFVVVVVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZnd3d3d3d4iIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d2ZmZoiIiIiIiHd3d3d3d3d3d2ZmZnd3d2ZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiJmZmZmZmZmZmZmZmZmZmYiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d2ZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d3d3d4iIiIiIiIiIiJmZmYiIiJmZmYiIiIiIiIiIiIiIiJmZmZmZmZmZmXd3d3d3d3d3d3d3d5mZmYiIiHd3d3d3d2ZmZmZmZmZmZmZmZnd3d3d3d4iIiHd3d4iIiIiIiJmZmaqqqqqqqpmZmaqqqpmZmYiIiJmZmYiIiHd3d4iIiHd3d4iIiHd3d4iIiHd3d4iIiHd3d4iIiHd3d4iIiHd3d3d3d3d3d4iIiHd3d4iIiHd3d4iIiHd3d2ZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d2ZmZlVVVVVVVVVVVVVVVVVVVURERERERERERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzM0RERDMzM0RERERERGZmZoiIiHd3d2ZmZlVVVWZmZmZmZmZmZlVVVURERFVVVVVVVURERDMzMzMzM0RERERERERERERERDMzM0RERGZmZru7u8zMzJmZmXd3d4iIiIiIiIiIiIiIiHd3d3d3d2ZmZlVVVVVVVWZmZlVVVURERERERFVVVVVVVURERERERERERFVVVURERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERDMzM0RERERERERERERERDMzM0RERDMzM0RERFVVVURERERERDMzMzMzMzMzMzMzM0RERERERERERFVVVVVVVVVVVVVVVWZmZlVVVXd3d5mZmXd3d2ZmZlVVVVVVVVVVVWZmZlVVVVVVVWZmZnd3d3d3d2ZmZkRERFVVVXd3d4iIiGZmZnd3d3d3d2ZmZlVVVURERERERDMzMzMzMzMzMzMzMzMzM0RERERERERERERERFVVVURERFVVVURERFVVVVVVVWZmZlVVVVVVVURERFVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d2ZmZmZmZnd3d4iIiHd3d3d3d3d3d4iIiIiIiIiIiFVVVURERERERFVVVVVVVVVVVURERERERERERERERERERERERERERERERERERERERERERFVVVURERERERERERERERERERERERERERERERERERERERERERFVVVVVVVURERERERERERFVVVURERFVVVURERFVVVURERERERERERFVVVURERERERERERFVVVVVVVVVVVVVVVXd3d3d3d3d3d4iIiIiIiIiIiHd3d4iIiIiIiHd3d3d3d3d3d2ZmZnd3d3d3d4iIiIiIiJmZmZmZmYiIiIiIiJmZmaqqqpmZmYiIiHd3d2ZmZmZmZnd3d4iIiHd3d2ZmZnd3d4iIiIiIiJmZmZmZmaqqqru7u7u7u8zMzMzMzMzMzLu7u6qqqpmZmZmZmaqqqt3d3f///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7u7u7u7u7d3d3d3d3d3d3d3d3u7u7d3d3d3d3d3d3u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3MzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7vMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3MzMzMzMzMzMyqqqqqqqqZmZmZmZmIiIiIiIiIiIiZmZmZmZmIiIiZmZmqqqqqqqqqqqqZmZmIiIh3d3dVVVVVVVVEREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNEREQzMzMzMzNVVVVVVVVERERERERVVVUzMzNERERERERVVVVVVVVVVVVVVVVERERERERERERVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZVVVVmZmZmZmZ3d3dmZmZmZmZmZmZmZmZ3d3eIiIh3d3d3d3d3d3eIiIh3d3eIiIiIiIiIiIh3d3dmZmZmZmZmZmZVVVVVVVVVVVVERERERERERERVVVVVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZ3d3eIiIiIiIiIiIh3d3eIiIiIiIiIiIiIiIiIiIiIiIiZmZmIiIiZmZmIiIiIiIiIiIiqqqq7u7vMzMyqqqqZmZmZmZmIiIhVVVVVVVVVVVVmZmZ3d3dmZmZVVVVmZmaqqqrMzMyZmZl3d3d3d3dmZmZVVVWIiIiIiIiIiIhmZmZVVVUzMzNERERmZmaIiIh3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVV3d3eIiIh3d3d3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZ3d3eIiIiIiIhmZmZVVVVmZmZmZmZVVVVERERERERVVVVVVVVVVVVVVVVVVVVmZmaIiIiIiIiIiIiIiIhmZmZVVVVmZmZmZmZmZmZmZmZmZmZVVVVERERERERERERVVVV3d3eIiIh3d3dmZmZmZmZmZmZERERERERVVVVVVVVVVVVVVVVERERERERVVVVmZmZ3d3dmZmZ3d3d3d3eZmZmIiIh3d3eIiIh3d3dmZmZ3d3d3d3dmZmZmZmZ3d3dmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3eIiIiIiIh3d3dmZmZVVVVmZmZmZmZVVVVmZmZVVVVmZmZmZmZ3d3dmZmZmZmZ3d3dmZmZmZmZmZmZmZmZ3d3d3d3eIiIiZmZmIiIiIiIh3d3dmZmZmZmZmZmZ3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3d3d3eIiIiZmZmIiIh3d3dmZmZmZmZ3d3d3d3dmZmZmZmZVVVVmZmZmZmZmZmZmZmZ3d3d3d3dmZmZ3d3d3d3d3d3eIiIh3d3dmZmZVVVVmZmZVVVVERERERERERERERERERERVVVVVVVVVVVVmZmZ3d3dmZmZVVVVmZmaIiIiIiIh3d3dmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3dmZmZVVVVmZmZ3d3eIiIhmZmZmZmZVVVVVVVVERERVVVVERERERERVVVVERERVVVVVVVVmZmZVVVVmZmZVVVVVVVVERERmZmaIiIiIiIhmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVmZmZmZmaIiIiIiIh3d3d3d3eIiIh3d3dmZmZVVVVmZmZmZmZmZmZ3d3d3d3dmZmZ3d3eIiIh3d3d3d3d3d3dmZmZ3d3eIiIiIiIh3d3eIiIiIiIh3d3d3d3dVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVEREQzMzMzMzNVVVVmZmZmZmZmZmZVVVVERERERERVVVVVVVVERERVVVVEREREREREREREREREREQzMzNEREREREREREREREQzMzMzMzNERERERERVVVVVVVVVVVVVVVVVVVVERERERERVVVVERERERERERERERERERERVVVVmZmZmZmZmZmZERERVVVVVVVVERERVVVVVVVVmZmZVVVVmZmZVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVmZmZVVVVVVVV3d3d3d3d3d3dVVVVVVVVmZmZVVVVmZmZVVVVmZmZmZmZ3d3d3d3d3d3d3d3dmZmZ3d3d3d3dmZmZ3d3eIiIiIiIh3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZmZmZ3d3d3d3d3d3eIiIiIiIiIiIiZmZmIiIiZmZmZmZmZmZmZmZmIiIiIiIiIiIh3d3eIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIiZmZmZmZmIiIh3d3eIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3eIiIiIiIiIiIiIiIiZmZmZmZmZmZmZmZmIiIiZmZmIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZVVVVVVVVVVVVVVVVEREREREREREREREREREREREREREREREQzMzNERERVVVVVVVVVVVVERERVVVVVVVVVVVV3d3eIiIhmZmZVVVVmZmaIiIiIiIhmZmZ3d3d3d3dmZmZVVVVEREQzMzMzMzNEREREREREREREREQzMzNVVVWZmZm7u7uqqqqZmZmIiIh3d3d3d3eIiIiIiIh3d3dmZmZVVVVVVVVVVVVVVVVEREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNEREQzMzNEREREREREREQzMzNERERERERERERERERVVVVEREREREQzMzMzMzMzMzNERERERERVVVVVVVVERERERERERERVVVVVVVVmZmZ3d3dmZmZmZmZmZmZVVVVERERmZmZERERVVVV3d3d3d3d3d3dmZmZVVVVVVVV3d3eIiIh3d3dmZmZmZmZmZmZVVVVEREREREQzMzMzMzMzMzNEREQzMzNERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3eIiIiIiIh3d3dVVVVERERERERVVVVEREREREREREREREQzMzNERERERERERERERERERERERERERERERERERERVVVVEREREREREREQzMzNERERERERERERERERERERERERVVVVERERERERERERERERVVVVERERERERVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVV3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIh3d3d3d3d3d3d3d3eIiIiIiIiIiIiZmZmZmZmZmZmZmZmZmZmZmZmqqqqIiIh3d3dVVVVmZmZmZmZmZmZmZmZmZmZ3d3eIiIiIiIiIiIiZmZmqqqq7u7vMzMzMzMzMzMy7u7uZmZl3d3eZmZmqqqrd3d3u7u7////////////////////u7u7////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u7u7u7u7u3d3d3d3dzMzMzMzM3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3d3d3dzMzMzMzMzMzMu7u7zMzMzMzMzMzM3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u3d3d7u7u3d3d3d3d3d3d3d3dzMzMzMzMu7u7u7u7u7u7qqqqqqqqqqqqqqqqmZmZmZmZmZmZiIiId3d3d3d3d3d3ZmZmVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREREREREREVVVVREREREREREREVVVVd3d3ZmZmZmZmZmZmVVVVZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiId3d3ZmZmZmZmZmZmd3d3ZmZmVVVVVVVVVVVVREREVVVVREREREREVVVVVVVVREREVVVVVVVVd3d3ZmZmZmZmZmZmVVVVVVVVZmZmVVVVREREREREVVVVREREVVVVVVVVVVVVZmZmVVVVZmZmZmZmd3d3ZmZmZmZmZmZmZmZmiIiId3d3d3d3d3d3iIiIiIiId3d3iIiIiIiIiIiIiIiIiIiImZmZmZmZmZmZd3d3d3d3iIiImZmZqqqqqqqqqqqqqqqqiIiId3d3d3d3VVVVZmZmiIiIiIiId3d3VVVVVVVVZmZmmZmZqqqqqqqqd3d3d3d3ZmZmREREd3d3d3d3d3d3VVVVREREREREREREZmZmd3d3d3d3d3d3ZmZmZmZmZmZmVVVVVVVVZmZmd3d3iIiIiIiIZmZmd3d3d3d3ZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVZmZmmZmZmZmZZmZmVVVVVVVVZmZmZmZmVVVVREREREREREREVVVVREREd3d3iIiId3d3d3d3iIiIiIiIZmZmREREZmZmZmZmZmZmZmZmZmZmZmZmREREREREVVVVZmZmd3d3ZmZmVVVVZmZmZmZmZmZmREREVVVVVVVVZmZmVVVVVVVVREREVVVVVVVVZmZmd3d3d3d3d3d3iIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmd3d3ZmZmZmZmZmZmd3d3ZmZmZmZmZmZmVVVVZmZmiIiIiIiId3d3d3d3ZmZmVVVVZmZmVVVVVVVVZmZmZmZmd3d3ZmZmd3d3d3d3d3d3d3d3ZmZmZmZmZmZmVVVVd3d3mZmZmZmZiIiIiIiIiIiIiIiId3d3ZmZmZmZmd3d3ZmZmZmZmd3d3ZmZmZmZmd3d3d3d3d3d3iIiImZmZiIiIiIiId3d3d3d3ZmZmZmZmd3d3ZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3iIiIiIiIiIiId3d3d3d3ZmZmVVVVVVVVREREREREREREVVVVVVVVVVVVZmZmd3d3d3d3VVVVZmZmiIiIiIiId3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3ZmZmZmZmd3d3d3d3d3d3ZmZmVVVVZmZmVVVVVVVVREREREREREREREREVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVZmZmd3d3d3d3ZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3iIiIZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVZmZmVVVVZmZmd3d3d3d3d3d3ZmZmd3d3d3d3d3d3ZmZmd3d3d3d3iIiId3d3ZmZmZmZmZmZmZmZmVVVVZmZmZmZmVVVVVVVVREREVVVVREREREREREREREREVVVVREREVVVVZmZmREREREREVVVVZmZmiIiId3d3ZmZmREREREREREREREREVVVVREREVVVVREREREREREREREREMzMzREREVVVVREREMzMzMzMzIiIiMzMzVVVVZmZmVVVVREREREREMzMzREREREREREREREREREREREREREREREREREREVVVVZmZmZmZmVVVVREREVVVVVVVVVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVd3d3iIiId3d3VVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmd3d3iIiId3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3iIiImZmZiIiImZmZiIiImZmZiIiImZmZmZmZiIiIiIiIiIiIiIiIiIiId3d3iIiId3d3d3d3d3d3d3d3d3d3ZmZmVVVVZmZmZmZmZmZmVVVVZmZmd3d3d3d3d3d3d3d3iIiIiIiId3d3iIiIiIiIiIiImZmZiIiIiIiIiIiIiIiId3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiImZmZiIiImZmZmZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmVVVVZmZmVVVVVVVVVVVVZmZmZmZmZmZmd3d3VVVVVVVVd3d3d3d3d3d3iIiIZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiIqqqqqqqqqqqqiIiIVVVVREREIiIiMzMzREREREREVVVVREREMzMzMzMzd3d3u7u7u7u7qqqqmZmZiIiIiIiId3d3iIiIiIiId3d3ZmZmVVVVVVVVVVVVREREREREREREVVVVREREMzMzREREREREVVVVVVVVREREREREVVVVREREMzMzREREREREMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREREREREREREREMzMzMzMzREREMzMzREREVVVVREREREREREREREREREREREREREREVVVVVVVVVVVVZmZmd3d3ZmZmVVVVREREREREZmZmd3d3d3d3ZmZmZmZmVVVVZmZmd3d3ZmZmZmZmZmZmVVVVVVVVREREREREMzMzMzMzREREREREMzMzREREREREREREREREVVVVREREVVVVREREVVVVVVVVVVVVREREVVVVREREREREVVVVREREVVVVVVVVREREVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVZmZmZmZmd3d3d3d3d3d3ZmZmVVVVREREREREREREREREREREREREREREREREREREMzMzREREREREMzMzREREMzMzREREREREVVVVREREREREREREREREREREMzMzREREREREREREREREREREREREVVVVREREVVVVREREREREVVVVVVVVREREVVVVREREVVVVVVVVVVVVVVVVZmZmd3d3d3d3ZmZmd3d3iIiIiIiIiIiImZmZmZmZqqqqmZmZmZmZmZmZiIiIiIiIiIiIiIiId3d3iIiImZmZmZmZmZmZqqqqqqqqmZmZmZmZmZmZqqqqiIiId3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3iIiImZmZqqqqu7u7u7u7u7u7iIiId3d3iIiImZmZu7u73d3d////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3e7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3d3d3d3d3czMzMzMzMzMzN3d3d3d3d3d3d3d3d3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3czMzMzMzLu7u7u7u6qqqpmZmYiIiHd3d2ZmZlVVVVVVVURERERERDMzMzMzMzMzMzMzMzMzM0RERERERERERDMzM0RERERERERERERERFVVVURERERERERERFVVVWZmZlVVVVVVVWZmZlVVVVVVVWZmZmZmZnd3d4iIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZlVVVWZmZmZmZnd3d4iIiHd3d4iIiIiIiHd3d4iIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d2ZmZmZmZlVVVURERERERFVVVURERERERERERERERERERERERFVVVVVVVVVVVVVVVURERERERFVVVWZmZmZmZlVVVVVVVVVVVURERFVVVURERFVVVVVVVWZmZlVVVWZmZlVVVWZmZnd3d2ZmZoiIiIiIiGZmZlVVVWZmZmZmZnd3d3d3d3d3d2ZmZmZmZnd3d2ZmZnd3d3d3d4iIiHd3d3d3d4iIiKqqqpmZmYiIiHd3d3d3d3d3d5mZmZmZmYiIiHd3d4iIiIiIiIiIiHd3d2ZmZmZmZoiIiIiIiGZmZmZmZlVVVVVVVXd3d4iIiIiIiHd3d3d3d2ZmZmZmZnd3d2ZmZmZmZmZmZkRERERERERERFVVVXd3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZpmZmYiIiGZmZmZmZmZmZnd3d2ZmZkRERERERFVVVWZmZmZmZmZmZlVVVWZmZmZmZoiIiGZmZmZmZlVVVWZmZmZmZmZmZlVVVURERERERERERFVVVWZmZmZmZlVVVWZmZnd3d3d3d2ZmZlVVVWZmZlVVVWZmZnd3d2ZmZnd3d2ZmZlVVVVVVVWZmZmZmZlVVVVVVVWZmZmZmZmZmZmZmZkRERFVVVVVVVVVVVVVVVVVVVURERFVVVWZmZnd3d3d3d4iIiIiIiIiIiHd3d2ZmZmZmZmZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZlVVVXd3d3d3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZnd3d3d3d2ZmZnd3d2ZmZmZmZlVVVWZmZmZmZnd3d4iIiJmZmYiIiHd3d3d3d4iIiIiIiHd3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZnd3d3d3d4iIiIiIiHd3d4iIiHd3d2ZmZmZmZnd3d2ZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d4iIiIiIiIiIiIiIiIiIiGZmZmZmZlVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d2ZmZlVVVWZmZmZmZmZmZlVVVWZmZlVVVURERFVVVVVVVWZmZmZmZmZmZnd3d2ZmZmZmZmZmZnd3d3d3d2ZmZlVVVVVVVWZmZmZmZlVVVVVVVVVVVURERERERERERFVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVXd3d3d3d1VVVVVVVVVVVVVVVWZmZmZmZlVVVWZmZlVVVURERERERERERFVVVVVVVVVVVWZmZnd3d2ZmZmZmZlVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVWZmZlVVVWZmZnd3d3d3d2ZmZnd3d3d3d2ZmZmZmZkRERFVVVVVVVWZmZmZmZlVVVVVVVURERERERERERERERERERERERERERERERFVVVVVVVXd3d3d3d1VVVVVVVWZmZlVVVVVVVVVVVURERFVVVURERERERERERERERFVVVURERERERERERERERERERERERERERDMzMzMzMzMzM1VVVWZmZmZmZkRERERERERERERERDMzMzMzMzMzM0RERDMzM0RERERERERERERERERERFVVVVVVVURERERERERERERERERERFVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d3d3d3d3d2ZmZnd3d2ZmZnd3d3d3d3d3d2ZmZmZmZlVVVWZmZlVVVWZmZmZmZlVVVVVVVVVVVWZmZnd3d2ZmZlVVVVVVVWZmZmZmZmZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d4iIiIiIiIiIiIiIiJmZmYiIiJmZmYiIiIiIiJmZmZmZmZmZmZmZmYiIiIiIiIiIiHd3d4iIiHd3d3d3d2ZmZmZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiJmZmYiIiIiIiJmZmYiIiJmZmYiIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiJmZmYiIiJmZmYiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZnd3d2ZmZmZmZnd3d2ZmZmZmZmZmZnd3d3d3d2ZmZmZmZmZmZmZmZlVVVWZmZlVVVWZmZnd3d3d3d2ZmZmZmZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZoiIiIiIiKqqqqqqqpmZmWZmZlVVVURERDMzMzMzMzMzM0RERFVVVURERDMzM0RERJmZmbu7u7u7u7u7u5mZmYiIiIiIiHd3d3d3d4iIiGZmZlVVVVVVVURERFVVVVVVVURERERERFVVVURERERERERERERERERERFVVVURERERERERERERERDMzMzMzM0RERDMzMzMzM0RERERERDMzMzMzM0RERERERDMzM0RERDMzMzMzMzMzM0RERDMzM0RERERERERERERERERERERERERERDMzM0RERERERERERERERERERERERERERERERERERERERERERERERDMzM0RERGZmZnd3d3d3d0RERERERFVVVURERGZmZmZmZoiIiGZmZlVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVURERDMzM0RERDMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERERERFVVVVVVVURERERERERERERERERERERERFVVVURERFVVVURERFVVVURERFVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVURERERERERERERERERERERERERERDMzMzMzM0RERFVVVURERERERERERERERERERERERERERDMzM0RERERERERERERERDMzM0RERDMzM0RERERERERERFVVVVVVVURERFVVVVVVVVVVVVVVVURERFVVVVVVVVVVVURERFVVVVVVVVVVVWZmZmZmZnd3d3d3d3d3d4iIiJmZmYiIiJmZmZmZmZmZmZmZmZmZmZmZmaqqqpmZmYiIiJmZmZmZmZmZmaqqqqqqqqqqqqqqqqqqqpmZmaqqqqqqqqqqqqqqqnd3d3d3d2ZmZmZmZnd3d3d3d2ZmZmZmZnd3d3d3d4iIiJmZmaqqqru7u7u7u7u7u5mZmXd3d2ZmZmZmZpmZmbu7u+7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7////u7u7////u7u7////u7u7////u7u7////u7u7////////u7u7d3d3d3d3MzMzd3d3MzMzd3d3d3d3d3d3u7u7u7u7u7u7u7u7d3d3u7u7d3d3MzMzMzMzMzMy7u7vMzMzMzMzMzMzd3d3d3d3d3d3d3d3d3d3u7u7d3d3d3d3MzMy7u7uqqqqIiIiIiIh3d3dVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzNERERERERVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZ3d3d3d3dmZmZmZmZ3d3d3d3dmZmZmZmZ3d3dmZmZmZmZ3d3d3d3eIiIiIiIh3d3eIiIiIiIh3d3d3d3d3d3d3d3eIiIh3d3eIiIiIiIiIiIh3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3eIiIiZmZmIiIiZmZmIiIiZmZmIiIiIiIiIiIh3d3dmZmZmZmZVVVVVVVVVVVVVVVVERERVVVVERERERERERERVVVVERERVVVVVVVVVVVVVVVVERERERERERERVVVVERERERERERERVVVVVVVVmZmZVVVVVVVVmZmZVVVVmZmZVVVV3d3d3d3d3d3d3d3dmZmZ3d3eIiIh3d3eIiIiIiIhmZmZVVVVmZmZ3d3d3d3d3d3dmZmZmZmZmZmZVVVVVVVV3d3d3d3d3d3d3d3eIiIiZmZmqqqqIiIiIiIh3d3eIiIiqqqqZmZmZmZl3d3dmZmZ3d3eIiIh3d3dmZmZmZmZVVVV3d3d3d3dmZmZVVVVVVVVVVVVmZmZmZmZVVVVmZmZmZmZ3d3eIiIh3d3dVVVVmZmZ3d3dVVVVERERVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmaIiIh3d3dmZmZmZmZmZmZmZmZVVVVVVVVERERVVVVmZmZVVVVVVVVVVVVVVVVmZmZ3d3dmZmZmZmZmZmZVVVVmZmZmZmZVVVVERERERERVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZVVVVmZmZVVVVVVVVVVVVmZmZ3d3d3d3dVVVVERERVVVVVVVVmZmZVVVVVVVVERERVVVVmZmZmZmZ3d3eIiIiIiIiIiIiIiIh3d3d3d3dmZmZmZmZVVVVmZmZmZmZmZmZmZmZ3d3eIiIhmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVVVVVmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmaIiIiIiIh3d3dmZmZmZmaIiIiIiIiIiIh3d3d3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIh3d3d3d3dmZmZ3d3dmZmZ3d3d3d3dmZmZmZmZ3d3dmZmZmZmZVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZ3d3dmZmZVVVVmZmZmZmZVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZ3d3dmZmZ3d3d3d3d3d3dmZmZVVVVERERVVVVVVVVVVVVmZmZVVVVVVVVERERERERERERVVVVVVVVmZmZVVVVmZmZVVVVVVVV3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVERERVVVVERERERERERERVVVVmZmZmZmZmZmZVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZ3d3eIiIh3d3dmZmZERERVVVVVVVVVVVVmZmZVVVVERERERERERERERERERERERERERERERERERERVVVVVVVV3d3dmZmZVVVVVVVVERERERERERERVVVVERERERERERERVVVVEREQzMzNEREREREREREREREQzMzNEREREREREREQzMzNEREREREREREREREREREQzMzNEREREREREREQzMzNERERERERERERERERERERERERERERERERERERERERERERERERVVVVVVVVEREQzMzMzMzMzMzNERERERERVVVVVVVVERERERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZVVVVmZmZVVVVVVVVVVVVmZmZVVVVmZmZmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZmZmZ3d3d3d3d3d3eIiIiIiIiIiIiIiIiZmZmZmZmZmZmZmZmZmZmIiIiZmZmIiIiIiIiIiIh3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3eIiIh3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZmIiIiZmZmIiIiIiIiZmZmIiIiZmZmIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZmZmZmIiIiZmZmIiIiZmZmIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3eIiIhmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3eIiIiIiIiIiIhmZmZEREQzMzMzMzMzMzNVVVVVVVVVVVVERERERER3d3eqqqq7u7u7u7uZmZmZmZmIiIiIiIiIiIiZmZl3d3dmZmZVVVVERERVVVVERERVVVVVVVVmZmZVVVVVVVVERERERERERERERERERERVVVVEREREREREREQzMzNEREQzMzMzMzMzMzMzMzNEREQzMzNEREQzMzNEREQzMzMzMzNEREQzMzMzMzNEREQzMzNEREQzMzNEREREREREREREREREREQzMzMzMzNEREQzMzNEREQzMzNERERERERERERVVVVEREQzMzNEREQzMzNVVVVVVVVVVVVERERERERERERVVVVVVVVmZmZmZmZmZmZmZmZVVVVmZmZ3d3dmZmZmZmZVVVVEREREREQzMzMzMzNEREQzMzMzMzMzMzNEREREREREREQzMzNERERERERERERERERERERVVVVERERERERERERERERERERERERERERERERERERVVVVERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVEREQzMzMzMzNERERERERERERVVVVEREQzMzNERERERERERERVVVVERERVVVVVVVVEREQzMzNEREQzMzNERERVVVVEREREREQzMzNEREQzMzNERERERERERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZ3d3d3d3dmZmZ3d3eIiIiIiIiZmZmIiIiZmZmZmZmIiIiIiIiZmZmIiIiIiIiIiIiIiIiIiIiZmZmqqqqqqqqqqqqqqqqZmZmZmZmqqqq7u7u7u7uZmZl3d3dmZmZ3d3d3d3eIiIh3d3d3d3eIiIiIiIiqqqqqqqqqqqq7u7u7u7uZmZl3d3dmZmZmZmZmZmaZmZnMzMzu7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u3d3d3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u7u7u7u7u3d3d3d3d3d3dzMzMu7u7u7u7u7u7zMzMzMzMzMzMzMzM3d3d3d3d3d3dzMzMzMzMzMzMzMzMu7u7u7u7qqqqiIiId3d3d3d3d3d3VVVVVVVVVVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3iIiIiIiId3d3d3d3d3d3iIiId3d3d3d3d3d3iIiId3d3d3d3iIiIiIiId3d3iIiIiIiIiIiIiIiIiIiId3d3iIiIiIiIiIiId3d3d3d3iIiId3d3d3d3iIiId3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZmZmZmZmZiIiIiIiIiIiId3d3VVVVVVVVVVVVREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVREREREREREREVVVVREREREREREREREREREREREREVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiId3d3d3d3iIiIZmZmd3d3ZmZmVVVVZmZmZmZmd3d3d3d3d3d3ZmZmd3d3ZmZmVVVVREREd3d3mZmZd3d3d3d3iIiIqqqqqqqqiIiIiIiImZmZqqqqqqqqmZmZiIiId3d3d3d3iIiImZmZiIiIZmZmZmZmZmZmd3d3ZmZmVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmd3d3d3d3ZmZmREREREREVVVVVVVVVVVVZmZmd3d3ZmZmZmZmZmZmZmZmVVVVd3d3ZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmd3d3ZmZmVVVVZmZmZmZmZmZmZmZmZmZmREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVZmZmd3d3d3d3d3d3ZmZmZmZmZmZmd3d3iIiId3d3d3d3VVVVZmZmVVVVZmZmd3d3d3d3d3d3VVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3d3d3d3d3iIiId3d3d3d3ZmZmZmZmVVVVZmZmZmZmd3d3ZmZmd3d3iIiId3d3ZmZmZmZmZmZmd3d3iIiId3d3ZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3ZmZmd3d3ZmZmd3d3ZmZmd3d3iIiId3d3d3d3ZmZmZmZmZmZmd3d3ZmZmZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVZmZmZmZmZmZmd3d3d3d3VVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmREREVVVVREREZmZmZmZmZmZmd3d3d3d3ZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVREREVVVVREREREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVREREVVVVREREVVVVZmZmVVVVZmZmVVVVVVVVREREVVVVREREREREVVVVZmZmZmZmZmZmVVVVREREMzMzREREREREREREREREREREVVVVVVVVVVVVVVVVREREREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmiIiIiIiIZmZmZmZmREREREREVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREREREMzMzREREVVVVZmZmZmZmVVVVVVVVREREREREMzMzREREREREREREREREREREREREREREREREMzMzREREREREREREMzMzMzMzMzMzREREVVVVREREREREREREMzMzMzMzIiIiMzMzREREREREREREREREREREMzMzREREREREREREREREREREREREREREREREREREVVVVREREMzMzMzMzMzMzMzMzREREVVVVVVVVVVVVREREREREREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVREREREREREREVVVVVVVVZmZmZmZmVVVVZmZmVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVZmZmd3d3ZmZmd3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3iIiIiIiIiIiIiIiImZmZmZmZmZmZmZmZmZmZmZmZiIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3iIiId3d3iIiIiIiImZmZiIiIiIiImZmZiIiImZmZiIiImZmZmZmZiIiImZmZmZmZmZmZmZmZmZmZmZmZiIiIiIiIiIiIiIiId3d3iIiId3d3iIiIiIiIiIiIiIiIiIiIiIiImZmZiIiImZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3ZmZmd3d3iIiIiIiId3d3d3d3d3d3ZmZmZmZmVVVVZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVREREVVVVZmZmVVVVVVVVREREZmZmVVVVZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmREREREREREREMzMzMzMzREREVVVVREREREREREREREREiIiIu7u7u7u7qqqqmZmZiIiIiIiId3d3qqqqmZmZZmZmVVVVVVVVVVVVVVVVREREVVVVZmZmVVVVVVVVREREREREREREREREREREREREREREMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzMzMzREREMzMzMzMzREREREREREREMzMzREREREREREREMzMzREREREREMzMzREREMzMzMzMzMzMzMzMzREREREREREREREREREREREREMzMzMzMzMzMzREREREREREREREREMzMzREREVVVVZmZmVVVVVVVVVVVVd3d3ZmZmZmZmZmZmREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREMzMzREREMzMzREREREREREREVVVVREREREREMzMzREREREREREREREREREREREREVVVVREREVVVVVVVVREREREREREREVVVVVVVVVVVVREREVVVVVVVVVVVVREREREREMzMzREREREREMzMzMzMzREREREREREREREREREREMzMzREREREREREREMzMzREREREREREREREREMzMzREREREREVVVVREREREREMzMzREREMzMzREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVZmZmZmZmZmZmd3d3iIiIiIiId3d3d3d3d3d3iIiImZmZiIiIiIiIiIiIiIiId3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3iIiImZmZqqqqu7u7qqqqqqqqqqqqqqqqu7u7qqqqqqqqiIiId3d3d3d3iIiIiIiIiIiImZmZqqqqu7u7u7u7u7u7u7u7mZmZd3d3d3d3ZmZmd3d3iIiImZmZu7u77u7u////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzN3d3czMzMzMzLu7u8zMzMzMzLu7u7u7u7u7u6qqqqqqqqqqqpmZmZmZmaqqqqqqqqqqqru7u6qqqqqqqpmZmZmZmZmZmYiIiIiIiHd3d4iIiIiIiIiIiJmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmYiIiJmZmaqqqpmZmYiIiIiIiIiIiIiIiHd3d4iIiHd3d4iIiIiIiIiIiJmZmYiIiIiIiIiIiIiIiIiIiHd3d4iIiHd3d4iIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiJmZmYiIiJmZmZmZmZmZmaqqqpmZmZmZmYiIiHd3d3d3d3d3d2ZmZlVVVVVVVVVVVURERERERERERERERERERERERERERFVVVVVVVVVVVVVVVWZmZlVVVURERERERFVVVURERERERERERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d2ZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d2ZmZlVVVVVVVWZmZnd3d3d3d2ZmZnd3d4iIiHd3d4iIiHd3d5mZmaqqqoiIiHd3d3d3d3d3d3d3d5mZmaqqqpmZmXd3d4iIiHd3d1VVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZkRERERERFVVVWZmZmZmZlVVVWZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVWZmZmZmZlVVVVVVVVVVVWZmZnd3d3d3d2ZmZlVVVURERFVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVWZmZnd3d3d3d2ZmZnd3d3d3d2ZmZmZmZnd3d4iIiHd3d2ZmZlVVVWZmZnd3d3d3d2ZmZmZmZlVVVVVVVVVVVVVVVURERFVVVVVVVWZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiGZmZmZmZmZmZmZmZmZmZmZmZnd3d4iIiIiIiGZmZlVVVWZmZnd3d3d3d2ZmZnd3d2ZmZnd3d3d3d2ZmZmZmZmZmZlVVVURERFVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZnd3d3d3d3d3d2ZmZnd3d3d3d2ZmZnd3d2ZmZnd3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZlVVVWZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVWZmZnd3d3d3d1VVVWZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d2ZmZmZmZlVVVURERFVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVWZmZlVVVURERERERFVVVURERFVVVWZmZmZmZmZmZlVVVVVVVURERFVVVVVVVURERFVVVURERFVVVVVVVVVVVVVVVWZmZlVVVVVVVURERERERFVVVWZmZlVVVVVVVURERDMzM0RERERERERERFVVVURERERERERERERERFVVVURERERERERERFVVVVVVVVVVVWZmZlVVVWZmZnd3d4iIiHd3d2ZmZkRERERERERERFVVVURERFVVVVVVVURERERERERERERERDMzM0RERDMzMzMzM1VVVVVVVVVVVVVVVWZmZlVVVURERERERDMzMzMzM0RERERERERERERERERERERERERERDMzM0RERDMzMzMzMzMzMzMzMzMzM1VVVVVVVVVVVTMzMzMzMzMzMzMzMzMzM0RERERERFVVVURERDMzMzMzM0RERDMzMzMzMzMzM0RERDMzM0RERERERERERFVVVURERERERERERERERERERERERDMzM1VVVVVVVVVVVVVVVURERERERERERDMzMzMzMzMzM0RERDMzMzMzM0RERFVVVURERERERERERERERERERDMzMzMzM0RERFVVVVVVVVVVVURERERERERERERERERERERERERERERERERERERERERERERERFVVVVVVVWZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVWZmZmZmZmZmZlVVVWZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVWZmZnd3d3d3d3d3d3d3d3d3d3d3d5mZmYiIiIiIiIiIiJmZmYiIiJmZmYiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiHd3d4iIiIiIiHd3d3d3d3d3d4iIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiJmZmYiIiJmZmYiIiJmZmYiIiJmZmZmZmZmZmYiIiJmZmYiIiIiIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiJmZmYiIiJmZmZmZmYiIiJmZmZmZmZmZmZmZmYiIiHd3d2ZmZmZmZlVVVWZmZlVVVVVVVVVVVWZmZmZmZlVVVWZmZlVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZlVVVURERDMzM0RERDMzMzMzM0RERFVVVVVVVURERDMzM0RERFVVVaqqqszMzKqqqqqqqoiIiIiIiIiIiJmZmZmZmXd3d1VVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERFVVVURERERERERERERERERERERERERERDMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERDMzM0RERERERERERDMzM0RERDMzM0RERERERERERERERERERERERERERDMzMzMzM0RERDMzM0RERERERERERERERFVVVURERDMzMzMzMzMzMzMzM0RERERERDMzMzMzMzMzM1VVVVVVVWZmZlVVVVVVVXd3d3d3d3d3d2ZmZlVVVURERERERERERDMzMzMzMzMzM0RERERERERERERERDMzMzMzMzMzM0RERERERERERERERERERERERERERERERDMzM0RERDMzM0RERERERERERERERERERERERFVVVURERERERERERFVVVURERERERERERERERDMzMzMzM0RERERERERERDMzM0RERERERERERERERERERERERERERERERERERERERDMzM0RERERERERERERERDMzM0RERERERERERERERDMzM0RERDMzM0RERERERFVVVURERFVVVVVVVURERFVVVURERFVVVURERFVVVVVVVVVVVWZmZnd3d4iIiIiIiIiIiHd3d4iIiHd3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZoiIiJmZmaqqqru7u6qqqqqqqqqqqru7u6qqqru7u6qqqpmZmYiIiIiIiJmZmZmZmaqqqru7u8zMzLu7u7u7u6qqqnd3d2ZmZmZmZnd3d3d3d5mZmbu7u93d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3MzMzMzMzMzMyqqqq7u7u7u7vMzMzMzMy7u7u7u7uqqqqqqqqZmZmZmZmZmZmZmZmZmZmZmZmqqqq7u7u7u7vMzMzMzMzMzMzMzMzd3d3MzMzMzMzMzMy7u7u7u7u7u7u7u7uqqqqqqqq7u7uqqqqqqqq7u7uqqqqqqqqqqqqqqqqqqqqZmZmqqqqZmZmZmZmZmZmZmZmZmZmIiIiIiIiIiIiZmZmIiIiZmZmqqqqZmZmZmZmZmZmIiIh3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3eIiIiIiIiIiIh3d3eIiIiIiIiIiIiIiIiIiIiIiIiZmZmZmZmZmZmZmZmZmZmIiIiZmZmIiIiIiIh3d3d3d3dmZmZVVVVmZmZVVVVmZmZVVVVVVVVERERVVVVERERERERVVVVVVVVERERVVVVERERVVVVVVVVERERVVVVERERVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVEREREREQzMzNERERERERVVVVVVVVmZmZmZmZmZmZmZmZ3d3eIiIiIiIiIiIh3d3dVVVVVVVVVVVV3d3d3d3eIiIiIiIhmZmZmZmZmZmZVVVV3d3eIiIiIiIh3d3dmZmZmZmZ3d3eZmZmqqqqZmZmIiIh3d3dmZmZVVVVVVVVVVVVERERERERVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZ3d3dmZmZ3d3dmZmZ3d3dmZmZmZmZVVVVERERVVVVVVVVVVVVERERVVVVmZmZ3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVERERVVVVVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3dmZmZmZmZmZmZ3d3dmZmZmZmZmZmZVVVVVVVVVVVVERERERERVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3eIiIh3d3dmZmZmZmZmZmZVVVVVVVV3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3eIiIh3d3dmZmZ3d3dmZmZ3d3d3d3dmZmZERERVVVVERERVVVVERERVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3eIiIhmZmZmZmZ3d3d3d3dmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZ3d3dmZmZmZmZ3d3dmZmZmZmZ3d3d3d3dmZmZ3d3d3d3d3d3d3d3dmZmZVVVVmZmZVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZmZmZVVVVERERVVVVmZmZmZmZmZmZVVVVmZmZmZmZVVVVmZmZVVVVVVVVmZmZ3d3d3d3d3d3dmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVmZmZ3d3dmZmZmZmZVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVERERERERERERmZmZmZmZmZmZVVVVVVVVVVVVERERVVVVERERERERERERERERERERVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVEREREREQzMzMzMzNERERERERERERERERERERERERERERERERVVVVERERERERVVVVVVVVmZmZVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVERERERERERERERERERERERERERERVVVVEREREREREREQzMzNEREQzMzNVVVVVVVVVVVVVVVVVVVVVVVVEREQzMzMzMzMzMzMzMzNERERVVVVEREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNVVVVEREREREREREREREREREREREQzMzNEREREREREREREREREREREREQzMzMzMzMzMzMzMzMzMzNEREQzMzNEREREREREREREREREREREREREREQzMzMzMzMzMzNERERVVVVVVVVVVVVEREREREQzMzMzMzNEREQzMzMzMzMzMzNERERERERVVVVEREREREREREREREQzMzMzMzMzMzNERERERERERERVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERVVVVVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3d3d3eIiIiIiIiIiIiZmZmIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3eIiIh3d3eIiIh3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZmZmZmIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZmZmZmZmZmZmZmIiIiIiIiZmZmIiIiZmZmIiIiIiIiIiIiIiIiIiIh3d3eIiIh3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZmZmZmIiIiIiIh3d3d3d3dmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZ3d3d3d3dmZmZVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZVVVVVVVVVVVVERERmZmZmZmZVVVVEREREREQzMzMzMzMzMzNERERVVVVVVVVERERERERERERERESIiIi7u7vMzMyqqqqIiIiIiIiIiIh3d3eZmZmIiIhmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZERERERERVVVVVVVVVVVVERERVVVVVVVVEREQiIiIzMzNEREQzMzMiIiIzMzMzMzMzMzMzMzNERERERERVVVVEREREREQzMzNEREQzMzMzMzNEREREREREREREREQzMzNEREREREREREREREREREQzMzNERERERERERERVVVVVVVVVVVVERERVVVVEREREREQzMzMzMzNERERVVVUzMzMzMzMzMzNERERVVVVVVVVVVVVVVVVVVVV3d3d3d3d3d3d3d3dmZmZVVVVEREQzMzMzMzMzMzNEREQzMzNEREQzMzNEREQzMzMzMzMzMzNEREREREREREREREREREREREQzMzNEREREREQzMzMzMzNEREQzMzMzMzNEREREREREREREREREREREREREREREREREREREREREREQzMzMzMzNEREQzMzNEREREREREREREREREREQzMzNEREREREREREREREQzMzNEREREREREREQzMzNEREQzMzNEREREREQzMzNEREQzMzNEREREREQzMzNERERERERVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVERERERERERERVVVVVVVV3d3eIiIiIiIiZmZmIiIiIiIh3d3dmZmZ3d3d3d3eIiIiIiIiIiIiIiIh3d3eIiIiIiIh3d3eIiIh3d3d3d3dmZmZ3d3d3d3eZmZmqqqqqqqq7u7uqqqq7u7u7u7uqqqq7u7uqqqqqqqqZmZmZmZmqqqqqqqq7u7u7u7vMzMy7u7uZmZmIiIhmZmZVVVV3d3d3d3eZmZmqqqq7u7vu7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////7u7u////7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3dzMzM3d3d3d3dzMzMzMzMu7u7mZmZmZmZmZmZmZmZmZmZmZmZd3d3iIiId3d3iIiImZmZmZmZqqqqu7u7zMzMzMzM3d3d3d3d3d3d3d3d3d3d7u7u3d3d3d3d3d3d3d3dzMzMzMzMu7u7u7u7u7u7u7u7u7u7qqqqqqqqu7u7qqqqqqqqu7u7qqqqu7u7qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqmZmZmZmZmZmZiIiIiIiIiIiId3d3d3d3ZmZmd3d3ZmZmZmZmd3d3d3d3d3d3d3d3iIiImZmZiIiImZmZiIiImZmZiIiImZmZmZmZiIiImZmZmZmZiIiIiIiId3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmREREREREREREVVVVVVVVREREREREREREREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVREREREREREREREREMzMzMzMzMzMzMzMzREREVVVVZmZmZmZmZmZmiIiId3d3ZmZmd3d3iIiId3d3ZmZmZmZmZmZmd3d3iIiImZmZiIiId3d3d3d3ZmZmVVVVREREZmZmiIiImZmZiIiIZmZmVVVVZmZmiIiIiIiId3d3ZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVREREREREVVVVVVVVVVVVREREVVVVREREVVVVVVVVREREREREVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmREREVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3ZmZmZmZmVVVVREREVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmVVVVVVVVREREVVVVVVVVZmZmZmZmd3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3ZmZmZmZmZmZmVVVVVVVVVVVVZmZmREREVVVVVVVVZmZmd3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3ZmZmVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3ZmZmZmZmd3d3iIiId3d3d3d3d3d3ZmZmd3d3iIiIZmZmVVVVREREREREREREVVVVREREVVVVVVVVZmZmZmZmVVVVZmZmd3d3iIiIiIiIZmZmZmZmd3d3iIiIZmZmZmZmZmZmd3d3d3d3ZmZmVVVVZmZmd3d3ZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmVVVVVVVVZmZmREREREREREREREREVVVVZmZmZmZmZmZmVVVVREREVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVREREREREd3d3iIiId3d3d3d3ZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmVVVVZmZmVVVVVVVVVVVVZmZmZmZmd3d3ZmZmZmZmd3d3ZmZmREREREREVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVREREREREREREREREREREREREREREREREVVVVREREREREVVVVZmZmd3d3VVVVVVVVZmZmZmZmVVVVREREREREMzMzREREREREREREVVVVVVVVREREREREREREREREVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmVVVVVVVVREREREREVVVVREREREREMzMzREREMzMzMzMzREREVVVVVVVVREREREREREREMzMzREREVVVVVVVVREREVVVVVVVVVVVVREREREREMzMzMzMzMzMzREREREREREREREREREREMzMzMzMzMzMzIiIiMzMzMzMzREREREREVVVVREREREREREREREREREREMzMzREREREREMzMzREREREREMzMzREREREREREREMzMzREREMzMzMzMzREREREREVVVVREREMzMzREREMzMzMzMzMzMzREREMzMzREREREREVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREVVVVREREREREREREREREMzMzMzMzMzMzMzMzREREREREVVVVREREREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREVVVVVVVVVVVVREREREREREREREREREREREREREREREREVVVVREREMzMzMzMzMzMzMzMzREREREREMzMzREREMzMzREREREREREREREREVVVVREREVVVVZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3iIiIiIiId3d3d3d3iIiId3d3iIiId3d3d3d3ZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVVVVVREREVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3iIiId3d3iIiIiIiImZmZiIiIiIiIiIiImZmZiIiImZmZmZmZmZmZmZmZiIiIiIiIiIiIiIiIiIiIiIiId3d3iIiId3d3d3d3d3d3d3d3iIiId3d3iIiId3d3iIiIiIiIiIiId3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiId3d3iIiIiIiIiIiIiIiImZmZiIiImZmZmZmZmZmZmZmZmZmZiIiIiIiIiIiIiIiId3d3iIiIiIiIiIiIiIiId3d3iIiImZmZiIiImZmZiIiId3d3d3d3ZmZmd3d3d3d3d3d3ZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmREREVVVVREREVVVVVVVVVVVVVVVVREREREREMzMzMzMzREREREREREREVVVVREREREREREREREREVVVVu7u7zMzMu7u7mZmZiIiId3d3d3d3iIiIiIiIZmZmZmZmVVVVVVVVZmZmVVVVREREZmZmd3d3VVVVREREREREREREREREVVVVVVVVZmZmREREMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREMzMzMzMzREREREREVVVVVVVVREREREREREREREREREREREREREREREREMzMzREREREREVVVVVVVVVVVVVVVVREREREREREREREREREREVVVVREREREREMzMzMzMzREREVVVVVVVVZmZmVVVVREREZmZmd3d3d3d3d3d3ZmZmVVVVREREREREMzMzMzMzMzMzMzMzREREREREREREMzMzMzMzMzMzREREMzMzREREREREREREREREREREMzMzMzMzREREMzMzMzMzREREREREREREREREREREMzMzREREREREREREREREREREREREREREMzMzREREMzMzREREMzMzREREREREREREREREREREMzMzREREMzMzREREREREREREMzMzREREREREMzMzREREMzMzREREMzMzMzMzREREREREREREREREREREMzMzREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmiIiImZmZmZmZiIiImZmZiIiId3d3iIiId3d3d3d3iIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3iIiImZmZqqqqu7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqu7u7qqqqu7u7u7u7u7u7zMzMzMzMqqqqiIiIZmZmZmZmVVVVd3d3iIiIqqqqu7u73d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////+7u7u7u7t3d3d3d3e7u7t3d3d3d3czMzN3d3czMzLu7u7u7u6qqqoiIiIiIiIiIiIiIiHd3d3d3d3d3d4iIiJmZmaqqqru7u8zMzMzMzN3d3e7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3bu7u7u7u8zMzLu7u7u7u6qqqru7u6qqqru7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqqqqqqqqqqqqqpmZmZmZmXd3d4iIiHd3d3d3d3d3d2ZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiIiIiIiIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZlVVVVVVVURERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVWZmZlVVVVVVVVVVVWZmZlVVVURERERERERERDMzMzMzMzMzM0RERERERERERERERERERERERDMzMzMzM0RERDMzM0RERERERERERFVVVURERFVVVWZmZoiIiHd3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d4iIiIiIiIiIiJmZmYiIiGZmZlVVVVVVVVVVVWZmZnd3d3d3d3d3d2ZmZmZmZmZmZnd3d3d3d2ZmZlVVVVVVVURERFVVVURERFVVVVVVVWZmZlVVVURERERERERERERERERERFVVVURERERERERERERERERERERERERERFVVVVVVVWZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZnd3d2ZmZlVVVVVVVURERFVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d2ZmZmZmZlVVVURERFVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVWZmZmZmZlVVVVVVVURERERERERERFVVVWZmZmZmZnd3d4iIiHd3d3d3d3d3d2ZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZlVVVWZmZlVVVVVVVVVVVWZmZmZmZlVVVVVVVURERGZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVXd3d3d3d3d3d3d3d2ZmZmZmZnd3d3d3d3d3d3d3d2ZmZlVVVVVVVVVVVURERFVVVWZmZmZmZlVVVURERERERFVVVWZmZnd3d4iIiIiIiIiIiHd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZnd3d3d3d3d3d2ZmZmZmZnd3d3d3d3d3d3d3d3d3d2ZmZlVVVWZmZlVVVWZmZlVVVVVVVURERERERERERGZmZnd3d2ZmZlVVVURERERERERERFVVVURERERERERERFVVVURERFVVVURERERERERERFVVVXd3d4iIiHd3d2ZmZlVVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVURERFVVVWZmZnd3d3d3d2ZmZmZmZlVVVURERERERERERFVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVWZmZmZmZmZmZlVVVURERFVVVURERERERERERERERERERFVVVURERFVVVVVVVURERFVVVVVVVWZmZlVVVWZmZlVVVVVVVVVVVTMzMzMzMzMzMzMzM0RERERERERERFVVVURERFVVVVVVVURERERERERERFVVVURERERERFVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERERERFVVVURERERERERERFVVVVVVVVVVVURERERERERERERERERERFVVVURERFVVVURERERERERERDMzM0RERERERERERERERERERERERERERDMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERDMzM0RERFVVVURERDMzM0RERERERDMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERDMzMzMzMzMzMzMzM0RERERERERERDMzM0RERDMzMzMzM0RERERERDMzMzMzM0RERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERDMzM0RERDMzMzMzMzMzMzMzM0RERERERDMzM0RERERERDMzMzMzMyIiIjMzMzMzMzMzMzMzM1VVVVVVVURERERERFVVVTMzM0RERDMzMzMzM0RERDMzM0RERERERERERDMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzM0RERERERDMzM0RERDMzMzMzM0RERDMzM0RERERERERERERERERERFVVVURERFVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d4iIiHd3d4iIiIiIiJmZmYiIiIiIiHd3d3d3d3d3d3d3d2ZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d4iIiIiIiIiIiJmZmYiIiJmZmZmZmZmZmZmZmZmZmYiIiJmZmZmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiHd3d3d3d3d3d3d3d3d3d4iIiHd3d4iIiHd3d3d3d3d3d3d3d4iIiHd3d4iIiIiIiIiIiIiIiIiIiJmZmZmZmZmZmYiIiIiIiJmZmYiIiIiIiIiIiJmZmYiIiIiIiIiIiJmZmZmZmYiIiIiIiGZmZmZmZlVVVWZmZmZmZnd3d3d3d3d3d2ZmZnd3d3d3d2ZmZmZmZmZmZnd3d3d3d2ZmZmZmZmZmZmZmZlVVVURERFVVVWZmZnd3d2ZmZlVVVTMzM0RERERERERERERERERERDMzM1VVVVVVVVVVVVVVVURERERERIiIiLu7u8zMzKqqqoiIiHd3d4iIiIiIiIiIiHd3d1VVVWZmZlVVVVVVVVVVVVVVVVVVVWZmZlVVVURERDMzM0RERFVVVVVVVWZmZkRERERERDMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERDMzM0RERERERERERERERERERERERDMzM0RERERERERERERERERERERERGZmZmZmZmZmZlVVVURERFVVVURERDMzM0RERFVVVVVVVVVVVTMzMzMzMzMzMzMzM1VVVVVVVVVVVVVVVVVVVURERGZmZnd3d2ZmZnd3d1VVVURERERERERERERERERERDMzM0RERERERDMzM0RERERERERERERERFVVVURERERERERERERERERERERERDMzMzMzM0RERERERDMzM0RERERERDMzM0RERDMzM0RERERERERERERERERERDMzM0RERDMzMzMzMzMzM0RERDMzM0RERERERERERERERDMzM0RERDMzM0RERERERERERERERERERFVVVURERERERDMzM0RERDMzM0RERDMzM0RERERERERERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVXd3d5mZmaqqqoiIiIiIiIiIiHd3d3d3d4iIiHd3d3d3d4iIiIiIiIiIiHd3d4iIiHd3d3d3d3d3d3d3d2ZmZmZmZnd3d4iIiJmZmZmZmaqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqru7u7u7u7u7u7u7u8zMzMzMzKqqqoiIiHd3d2ZmZmZmZmZmZoiIiKqqqru7u93d3e7u7u7u7v///////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////u7u7u7u7d3d3d3d3d3d3d3d3MzMzMzMzMzMy7u7uqqqqZmZmIiIh3d3d3d3eIiIiIiIiqqqqZmZmZmZmqqqq7u7vMzMzu7u7d3d3u7u7d3d3u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3MzMzMzMzd3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7uqqqqqqqqZmZmIiIiIiIiIiIh3d3d3d3d3d3eIiIh3d3d3d3dmZmZ3d3eIiIiIiIiZmZmIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3dmZmZ3d3dmZmZVVVVmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVERERERERVVVVERERVVVVERERERERVVVVERERERERVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZEREREREREREQzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNERERERERVVVVVVVVVVVVVVVVERERERERVVVV3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmaIiIiZmZl3d3dmZmZERERVVVVmZmZmZmZmZmZVVVVmZmZ3d3dmZmZmZmZVVVVVVVVmZmZVVVVVVVVVVVVERERVVVVmZmZVVVVVVVVVVVVVVVVERERERERERERERERVVVVERERVVVUzMzNERERERERERERERERERERVVVVmZmZmZmZ3d3dmZmZ3d3d3d3eIiIh3d3dmZmZ3d3dmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZERERERERVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZVVVVERERERERERERVVVVERERVVVVmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVERERVVVV3d3d3d3dmZmZVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZVVVVVVVVVVVVmZmZ3d3d3d3dVVVVVVVVVVVVmZmZ3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZERERERERVVVVVVVV3d3d3d3d3d3eIiIh3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVERERVVVVVVVVmZmZ3d3dmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZVVVVmZmZVVVVVVVVVVVVVVVVERERERERERERERERmZmZmZmZVVVUzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzNERERVVVV3d3d3d3d3d3dVVVVERERERERVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVmZmZmZmZ3d3dVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVERERERERERERERERVVVVmZmZmZmZERERERERVVVVERERERERERERERERERERERERERERERERVVVVVVVVERERERERVVVVERERVVVVmZmZmZmZmZmZVVVVEREQzMzMzMzMzMzNERERERERERERVVVVERERVVVVVVVVEREQzMzMzMzNERERERERVVVVmZmZVVVVVVVVEREQzMzNEREQzMzNERERERERERERERERERERERERVVVVERERERERERERERERVVVVERERVVVVERERVVVVVVVVVVVVERERERERERERERERERERERERERERERERVVVVVVVVEREREREREREREREREREQzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzNEREREREREREQzMzMzMzMzMzMzMzNEREQzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzNVVVVVVVVVVVVEREREREQzMzNEREREREQzMzNEREREREREREQzMzNEREREREQzMzMzMzMzMzNEREREREREREREREQzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNEREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNEREREREREREQzMzNEREQzMzMzMzMzMzNEREQzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNEREREREQzMzMzMzMzMzNEREQzMzNEREQzMzNERERVVVVERERERERERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3dmZmZ3d3eIiIh3d3d3d3eIiIiIiIh3d3eIiIiIiIh3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3eIiIiIiIiIiIiIiIiZmZmZmZmIiIiZmZmZmZmIiIiIiIiIiIiIiIiZmZmIiIiZmZmZmZmIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3eIiIh3d3d3d3d3d3dmZmZ3d3dmZmZ3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIiZmZmIiIiZmZmIiIiZmZmZmZmIiIiZmZmIiIiZmZmZmZmZmZmIiIh3d3d3d3dmZmZVVVVVVVVmZmZmZmZ3d3d3d3dmZmZVVVVmZmZmZmZmZmZVVVV3d3d3d3dmZmZVVVVVVVVmZmZVVVVVVVVmZmZmZmZmZmZmZmZVVVVEREREREQzMzNEREREREREREQzMzNERERVVVVERERVVVVERERERER3d3e7u7vMzMyqqqqIiIhmZmZ3d3eIiIiZmZmIiIhmZmZVVVVmZmZmZmZVVVVVVVVmZmZmZmZVVVVEREQzMzNERERERERVVVVEREREREREREREREQzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzNEREQzMzNEREQzMzNEREQzMzNEREQzMzNEREREREREREQzMzNERERVVVVEREQzMzNEREREREQzMzNERERERERVVVVmZmZmZmZmZmZVVVVERERERERERERERERERERmZmZmZmZEREQzMzMzMzMzMzNERERVVVVVVVVVVVVmZmZmZmZVVVVVVVVmZmZmZmZVVVVVVVVVVVVERERERERERERERERERERERERERERERERERERERERVVVVVVVVVVVVEREREREREREREREQzMzMzMzMzMzNEREQzMzMzMzNEREREREREREREREREREREREREREREREREREQzMzNEREREREREREQzMzMzMzMzMzNEREQzMzNEREREREQzMzNEREREREREREREREREREREREQzMzNEREREREREREREREREREREREREREREREQzMzNERERVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZmZmaIiIiZmZmZmZmIiIiIiIiIiIh3d3eIiIiIiIh3d3eIiIiIiIiIiIiIiIh3d3d3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3eIiIiIiIiZmZmqqqqZmZmZmZmZmZmqqqqqqqq7u7u7u7u7u7vMzMzMzMy7u7uqqqqIiIhmZmZmZmZmZmZ3d3eIiIiZmZm7u7vMzMzu7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7uzMzMzMzMu7u7zMzMzMzMu7u7u7u7qqqqmZmZd3d3d3d3d3d3iIiImZmZqqqqu7u7zMzMzMzMzMzM3d3d7u7u7u7u7u7u7u7u3d3d7u7u7u7u3d3d3d3d7u7u3d3d3d3d3d3d3d3dzMzMzMzM3d3dzMzM3d3dzMzM3d3d3d3dzMzM3d3dzMzMzMzM3d3dzMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7qqqqqqqqqqqqmZmZqqqqqqqqmZmZmZmZiIiImZmZiIiIiIiIiIiIiIiIiIiId3d3iIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVREREVVVVREREVVVVREREVVVVREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVZmZmVVVVREREVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmZmZmd3d3d3d3d3d3ZmZmVVVVVVVVVVVVREREVVVVMzMzMzMzMzMzMzMzREREREREVVVVREREMzMzREREREREMzMzMzMzMzMzREREREREREREVVVVVVVVVVVVREREREREZmZmd3d3ZmZmVVVVZmZmVVVVZmZmZmZmVVVVZmZmVVVVZmZmZmZmZmZmiIiIiIiId3d3ZmZmREREVVVVZmZmVVVVREREVVVVZmZmZmZmVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVd3d3d3d3VVVVREREREREREREREREREREREREVVVVREREVVVVVVVVREREREREREREREREREREVVVVVVVVVVVVZmZmZmZmd3d3d3d3iIiId3d3d3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmd3d3ZmZmVVVVREREVVVVREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVREREREREREREREREVVVVVVVVVVVVZmZmZmZmd3d3d3d3iIiId3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVZmZmd3d3d3d3VVVVVVVVVVVVZmZmd3d3ZmZmd3d3d3d3ZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVREREVVVVREREVVVVd3d3d3d3ZmZmd3d3d3d3ZmZmZmZmVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmREREVVVVVVVVZmZmZmZmZmZmVVVVZmZmVVVVZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREZmZmZmZmVVVVMzMzMzMzMzMzMzMzREREMzMzREREMzMzMzMzREREMzMzMzMzMzMzREREVVVVVVVVd3d3ZmZmZmZmVVVVREREREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREVVVVZmZmd3d3VVVVREREVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmVVVVREREMzMzMzMzREREVVVVVVVVZmZmVVVVREREREREREREREREREREREREREREREREREREREREREREVVVVREREREREREREREREREREVVVVZmZmZmZmVVVVREREMzMzMzMzREREREREREREREREVVVVREREVVVVVVVVREREMzMzMzMzIiIiREREVVVVZmZmZmZmREREMzMzREREMzMzMzMzREREREREREREREREVVVVREREREREREREREREMzMzREREMzMzREREREREVVVVVVVVVVVVREREREREREREREREREREVVVVVVVVVVVVREREMzMzREREREREMzMzREREMzMzMzMzVVVVREREREREREREMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREMzMzVVVVd3d3d3d3REREMzMzREREMzMzREREREREREREREREREREREREMzMzMzMzMzMzREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzREREMzMzMzMzMzMzREREREREMzMzREREMzMzREREREREREREMzMzMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3iIiId3d3iIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmd3d3ZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVd3d3d3d3iIiIiIiId3d3iIiImZmZiIiIiIiIiIiImZmZiIiImZmZiIiIiIiImZmZiIiIiIiIiIiImZmZiIiImZmZiIiImZmZiIiImZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3ZmZmZmZmd3d3iIiId3d3iIiIiIiIiIiIiIiIiIiIiIiId3d3iIiId3d3iIiIiIiIiIiIiIiId3d3iIiIiIiId3d3d3d3d3d3ZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmd3d3d3d3d3d3VVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVREREMzMzREREREREREREMzMzREREREREVVVVREREREREREREZmZmqqqqzMzMu7u7iIiIiIiId3d3iIiImZmZiIiIZmZmZmZmVVVVVVVVVVVVZmZmVVVVZmZmREREREREREREREREVVVVREREREREMzMzREREREREVVVVMzMzMzMzREREREREMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREREREREREREREREREMzMzMzMzMzMzREREREREVVVVREREVVVVVVVVVVVVVVVVREREVVVVREREREREVVVVZmZmVVVVMzMzMzMzMzMzREREREREREREVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREVVVVZmZmVVVVREREVVVVVVVVZmZmZmZmVVVVVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREREREREREREREREREREREREREREREREREMzMzREREMzMzREREREREREREMzMzREREREREMzMzREREREREREREREREREREMzMzREREMzMzREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVREREVVVVVVVVZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmiIiImZmZmZmZmZmZiIiIiIiId3d3iIiIiIiIiIiImZmZmZmZmZmZiIiId3d3d3d3d3d3ZmZmZmZmd3d3iIiId3d3iIiIiIiIiIiImZmZmZmZmZmZmZmZmZmZmZmZqqqqu7u7u7u7zMzMzMzMqqqqqqqqiIiId3d3ZmZmZmZmd3d3iIiImZmZqqqqzMzM3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////+7u7t3d3bu7u7u7u6qqqru7u7u7u6qqqqqqqqqqqpmZmZmZmYiIiJmZmaqqqru7u8zMzMzMzO7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqru7u6qqqqqqqqqqqqqqqqqqqpmZmaqqqpmZmaqqqpmZmZmZmZmZmZmZmYiIiIiIiIiIiIiIiHd3d4iIiHd3d2ZmZlVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVURERERERERERERERERERDMzMzMzM0RERERERERERERERERERERERERERERERERERFVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d2ZmZmZmZnd3d3d3d2ZmZmZmZlVVVURERERERERERERERERERERERERERERERERERERERFVVVVVVVURERERERERERERERERERERERDMzMzMzMzMzMzMzM0RERFVVVWZmZmZmZlVVVVVVVWZmZnd3d2ZmZlVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d3d3d3d3d2ZmZkRERERERERERERERDMzM0RERFVVVURERERERGZmZoiIiHd3d2ZmZlVVVWZmZmZmZmZmZlVVVVVVVURERFVVVVVVVURERERERERERERERFVVVURERFVVVWZmZkRERFVVVURERFVVVURERERERFVVVVVVVWZmZnd3d3d3d5mZmXd3d3d3d2ZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d3d3d3d3d2ZmZlVVVVVVVVVVVURERFVVVWZmZmZmZmZmZnd3d2ZmZmZmZlVVVWZmZmZmZmZmZkRERERERERERERERFVVVURERFVVVWZmZmZmZnd3d2ZmZmZmZnd3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZnd3d2ZmZnd3d2ZmZnd3d2ZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVWZmZlVVVURERFVVVVVVVXd3d2ZmZmZmZlVVVWZmZmZmZmZmZnd3d2ZmZnd3d2ZmZmZmZmZmZlVVVURERERERFVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d3d3d2ZmZlVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVURERFVVVWZmZmZmZlVVVURERDMzMzMzM0RERERERERERDMzMzMzM0RERFVVVVVVVTMzM0RERERERFVVVVVVVXd3d3d3d1VVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERFVVVWZmZmZmZlVVVURERFVVVURERFVVVURERFVVVVVVVURERFVVVVVVVVVVVVVVVURERERERDMzMzMzM0RERERERFVVVWZmZlVVVURERERERDMzMzMzMzMzM0RERERERERERDMzM0RERERERERERERERERERDMzM0RERERERFVVVVVVVWZmZlVVVURERDMzMzMzM0RERDMzM0RERERERERERFVVVURERERERERERDMzMzMzMzMzM0RERFVVVVVVVVVVVVVVVURERERERDMzM0RERDMzM0RERERERERERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVURERERERDMzMzMzM0RERFVVVURERDMzM0RERDMzM0RERDMzM0RERERERDMzM0RERERERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERERERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVURERFVVVURERERERGZmZnd3d1VVVURERERERDMzM0RERERERERERDMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVURERERERDMzMzMzM0RERERERERERERERDMzM0RERDMzMzMzMzMzMzMzM0RERERERDMzMyIiIjMzMzMzM0RERFVVVVVVVURERDMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERERERERERERERFVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d2ZmZmZmZmZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVURERFVVVURERERERFVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d2ZmZnd3d3d3d3d3d4iIiHd3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZnd3d2ZmZmZmZlVVVWZmZnd3d3d3d4iIiHd3d3d3d3d3d3d3d3d3d4iIiIiIiHd3d4iIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d2ZmZmZmZnd3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d2ZmZnd3d2ZmZnd3d4iIiJmZmaqqqoiIiHd3d3d3d2ZmZmZmZlVVVVVVVVVVVWZmZmZmZlVVVURERERERERERERERDMzMzMzM0RERERERDMzM0RERERERERERFVVVaqqqszMzMzMzJmZmZmZmYiIiIiIiJmZmYiIiGZmZmZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERDMzM1VVVVVVVURERERERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERDMzM0RERDMzM0RERERERERERERERERERERERDMzMzMzMzMzMzMzM0RERERERERERFVVVVVVVVVVVVVVVVVVVVVVVURERFVVVWZmZmZmZlVVVTMzMzMzMzMzMzMzM0RERGZmZmZmZlVVVWZmZlVVVVVVVURERFVVVVVVVVVVVWZmZlVVVURERERERERERERERFVVVVVVVURERFVVVVVVVWZmZmZmZnd3d2ZmZlVVVWZmZlVVVTMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERERERERERDMzM0RERERERERERERERFVVVVVVVURERFVVVURERDMzMzMzMzMzM0RERERERERERERERERERERERERERERERERERERERERERFVVVURERERERFVVVURERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZmZmZnd3d2ZmZnd3d2ZmZmZmZmZmZmZmZoiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiIiIiIiIiJmZmXd3d4iIiIiIiHd3d2ZmZnd3d2ZmZmZmZnd3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiJmZmaqqqru7u7u7u7u7u7u7u5mZmXd3d2ZmZmZmZmZmZnd3d5mZmZmZmaqqqru7u93d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d27u7vMzMzMzMzMzMy7u7vMzMy7u7u7u7u7u7u7u7vMzMzd3d3u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7u7u7u7u7d3d3d3d3d3d3d3d3MzMzd3d3d3d3MzMzd3d3MzMzMzMzMzMy7u7u7u7uqqqq7u7u7u7u7u7u7u7u7u7vMzMy7u7u7u7u7u7u7u7vMzMy7u7u7u7u7u7uqqqq7u7uqqqqZmZmZmZmZmZmIiIiIiIiIiIh3d3dmZmZVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVEREREREREREREREREREREREQzMzNERERERERERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZVVVVVVVVVVVVERERVVVVmZmZmZmZ3d3dmZmZ3d3eIiIh3d3dmZmZmZmZVVVVEREREREQzMzMzMzMzMzMzMzMzMzNERERVVVVERERVVVVVVVVERERERERVVVUzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzNERERVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZ3d3d3d3dVVVVVVVVVVVVVVVV3d3dmZmZmZmZVVVVVVVVEREQzMzMiIiJERERERERERERERER3d3eZmZmZmZmIiIhmZmZ3d3dmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVERERERERERERERERmZmZmZmZVVVVVVVVVVVVERERERERERERERERERERVVVVmZmZ3d3d3d3eIiIh3d3d3d3d3d3dmZmZmZmZ3d3eIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3eIiIh3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3d3d3dVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZmZmZmZmZ3d3d3d3dmZmZmZmZmZmZERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZ3d3d3d3dmZmZVVVV3d3dmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERVVVVmZmZVVVVERERVVVVVVVVmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVV3d3d3d3dmZmZEREREREQzMzMzMzNVVVVEREREREQzMzNERERERERmZmZEREQzMzNERERERERVVVV3d3dmZmZmZmZmZmZERERERERVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVERERERERERERERERERERERERmZmZmZmZVVVVVVVVVVVVERERERERERERERERERERERERERERERERERERVVVVEREQzMzMzMzNEREQzMzMzMzNVVVVmZmZVVVVEREQzMzMzMzNEREREREQzMzNEREREREQzMzNEREREREREREREREQzMzNERERERERERERERERVVVVVVVVVVVVEREREREQzMzNEREREREREREREREREREREREREREREREQzMzMiIiIiIiIzMzNERERVVVVVVVVVVVVEREREREQzMzNEREQzMzMzMzNEREREREREREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVVVVVEREQzMzMzMzMzMzNEREQzMzNEREREREQzMzNEREQzMzMzMzMzMzNEREREREQzMzMzMzNERERERERERERERERVVVVEREQzMzMzMzMzMzMzMzNEREREREREREREREREREQzMzNEREREREREREQzMzMzMzMiIiIzMzMzMzMzMzNERERVVVVERERERERmZmZmZmZEREQzMzMzMzNEREREREQzMzNEREREREQzMzMzMzMzMzMiIiIiIiIiIiIzMzNERERERERERERVVVVEREQzMzNEREQzMzMzMzNEREQzMzNEREQzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzMiIiIiIiIiIiIzMzNERERVVVVEREQzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzNERERERERERERERERERERERERVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVVVVVmZmZVVVVVVVVVVVVEREREREREREREREREREREREREREQzMzNERERERERERERERERVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dmZmaIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIh3d3eIiIh3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIh3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3eIiIh3d3eIiIh3d3d3d3eIiIiIiIiIiIh3d3eIiIh3d3d3d3dmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVmZmZmZmZ3d3d3d3eIiIiIiIh3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIiZmZmqqqqZmZmZmZmZmZl3d3dmZmZmZmZVVVVmZmZ3d3dmZmZERERERERVVVVVVVUzMzMzMzNEREREREREREQzMzMzMzMzMzMzMzNVVVWZmZnMzMzMzMyqqqqZmZmIiIiZmZmZmZmZmZl3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVEREREREREREREREQzMzNERERVVVVVVVVEREQzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzNEREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzNERERERERERERERERVVVVmZmZmZmZmZmZVVVVERERVVVVmZmZ3d3dVVVUzMzMzMzNERERERERVVVV3d3dmZmZmZmZmZmZVVVVVVVVERERERERmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVVERERERERERERVVVV3d3d3d3d3d3d3d3dmZmZVVVVEREQzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzNEREREREQzMzNERERERERVVVVVVVVVVVVVVVVEREREREREREREREQzMzNERERERERERERERERERERVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3eIiIh3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3eIiIh3d3eIiIh3d3eIiIiIiIiZmZmqqqqqqqqqqqqZmZmIiIhmZmZmZmZmZmZmZmZ3d3eZmZmqqqq7u7vMzMzMzMzd3d3u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u3d3d7u7u3d3d7u7u3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7zMzMzMzMzMzMzMzMzMzMzMzMu7u7zMzMu7u7u7u7u7u7qqqqqqqqqqqqmZmZiIiIiIiId3d3ZmZmZmZmVVVVVVVVREREVVVVREREVVVVVVVVVVVVVVVVREREREREVVVVREREVVVVREREREREVVVVREREREREREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3ZmZmZmZmVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVVVVVVVVVREREREREREREMzMzMzMzREREMzMzREREVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVZmZmVVVVVVVVZmZmVVVVVVVVZmZmiIiId3d3ZmZmVVVVZmZmZmZmVVVVVVVVREREREREVVVVZmZmd3d3ZmZmVVVVREREVVVVREREIiIiMzMzVVVVVVVVVVVVZmZmd3d3iIiId3d3ZmZmZmZmZmZmVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmREREREREVVVVVVVVVVVVREREREREVVVVVVVVZmZmZmZmZmZmd3d3d3d3iIiIiIiIiIiImZmZmZmZmZmZmZmZmZmZqqqqmZmZqqqqmZmZmZmZqqqqqqqqmZmZmZmZiIiId3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmZmZmVVVVREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3ZmZmZmZmd3d3ZmZmd3d3d3d3iIiId3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3iIiId3d3VVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmVVVVVVVVVVVVZmZmd3d3ZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVZmZmd3d3ZmZmZmZmZmZmd3d3ZmZmZmZmVVVVZmZmZmZmVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVd3d3d3d3ZmZmVVVVREREREREREREREREREREREREMzMzMzMzMzMzREREREREMzMzMzMzREREZmZmd3d3ZmZmZmZmVVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREREREREREREREVVVVZmZmVVVVVVVVREREVVVVREREVVVVREREVVVVREREREREREREREREVVVVREREREREREREMzMzMzMzREREVVVVZmZmVVVVREREREREMzMzREREREREREREREREMzMzREREMzMzREREREREREREREREREREMzMzREREVVVVREREVVVVVVVVREREMzMzMzMzREREREREREREREREREREREREREREREREMzMzIiIiMzMzMzMzMzMzVVVVVVVVVVVVVVVVREREMzMzMzMzREREREREMzMzREREMzMzREREREREMzMzREREMzMzMzMzREREMzMzREREMzMzREREZmZmVVVVREREREREMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREMzMzMzMzMzMzREREREREREREREREREREREREMzMzREREMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzREREREREREREREREd3d3iIiIZmZmREREMzMzREREMzMzREREMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzIiIiIiIiMzMzMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzVVVVZmZmVVVVREREVVVVVVVVREREVVVVVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVZmZmZmZmZmZmZmZmVVVVZmZmVVVVZmZmZmZmd3d3ZmZmZmZmZmZmVVVVREREVVVVVVVVREREREREREREREREREREREREREREREREREREVVVVREREREREMzMzREREREREREREREREVVVVVVVVZmZmVVVVZmZmVVVVZmZmZmZmd3d3d3d3iIiId3d3d3d3d3d3iIiIiIiId3d3iIiIiIiIiIiIiIiId3d3iIiId3d3iIiId3d3iIiId3d3iIiId3d3d3d3d3d3d3d3d3d3iIiId3d3iIiId3d3d3d3iIiId3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiId3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiImZmZiIiIiIiIiIiId3d3d3d3iIiId3d3d3d3ZmZmVVVVZmZmd3d3d3d3ZmZmVVVVZmZmVVVVREREMzMzMzMzREREREREMzMzIiIiMzMzMzMzREREVVVViIiIzMzMzMzMu7u7mZmZiIiImZmZqqqqmZmZZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVREREREREREREREREREREMzMzREREVVVVREREMzMzREREMzMzREREVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVVVVVVVVVZmZmVVVVVVVVVVVVREREZmZmZmZmZmZmVVVVREREMzMzMzMzREREVVVVd3d3ZmZmVVVVVVVVVVVVZmZmVVVVREREZmZmZmZmZmZmZmZmVVVVVVVVZmZmd3d3ZmZmZmZmREREREREREREVVVVVVVVd3d3iIiIiIiId3d3VVVVREREMzMzMzMzMzMzMzMzREREREREREREMzMzREREREREREREREREREREVVVVREREVVVVVVVVREREREREREREREREVVVVREREMzMzREREREREREREREREVVVVVVVVZmZmVVVVVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVZmZmREREREREVVVVZmZmVVVVVVVVZmZmiIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3iIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmZmZmd3d3ZmZmZmZmd3d3ZmZmiIiId3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3iIiIiIiImZmZmZmZqqqqmZmZiIiId3d3ZmZmVVVVVVVVZmZmd3d3iIiImZmZzMzM3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7v///////////////////+7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3d3d3e7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzN3d3czMzMzMzMzMzMzMzMzMzLu7u8zMzMzMzLu7u7u7u8zMzLu7u8zMzMzMzMzMzMzMzMzMzLu7u8zMzMzMzLu7u7u7u7u7u7u7u6qqqpmZmZmZmYiIiHd3d2ZmZlVVVVVVVURERFVVVURERERERERERERERERERERERERERFVVVURERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVXd3d3d3d2ZmZlVVVWZmZlVVVXd3d2ZmZnd3d3d3d2ZmZnd3d2ZmZmZmZlVVVURERERERERERDMzM0RERERERERERERERERERFVVVURERERERERERERERERERERERERERFVVVVVVVURERERERERERFVVVURERERERERERFVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVWZmZmZmZmZmZoiIiJmZmXd3d2ZmZlVVVWZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVWZmZnd3d1VVVURERFVVVWZmZkRERDMzM1VVVWZmZlVVVVVVVWZmZnd3d2ZmZmZmZmZmZlVVVVVVVVVVVURERERERERERFVVVWZmZmZmZlVVVWZmZmZmZlVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVWZmZnd3d3d3d4iIiIiIiJmZmZmZmaqqqszMzMzMzMzMzMzMzN3d3czMzMzMzLu7u7u7u7u7u8zMzLu7u7u7u8zMzLu7u7u7u6qqqqqqqpmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiGZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVURERFVVVWZmZlVVVWZmZmZmZlVVVWZmZmZmZmZmZlVVVWZmZmZmZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZnd3d3d3d3d3d3d3d2ZmZnd3d2ZmZnd3d2ZmZmZmZlVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVWZmZnd3d3d3d1VVVVVVVVVVVWZmZnd3d2ZmZmZmZmZmZlVVVVVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZnd3d3d3d1VVVVVVVWZmZlVVVVVVVWZmZmZmZlVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d2ZmZlVVVVVVVVVVVURERFVVVVVVVVVVVVVVVURERFVVVURERERERFVVVVVVVVVVVWZmZlVVVVVVVWZmZmZmZmZmZlVVVVVVVURERERERERERERERERERERERDMzMzMzMzMzMzMzM0RERDMzM0RERFVVVXd3d3d3d2ZmZlVVVURERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERFVVVWZmZlVVVVVVVURERFVVVURERFVVVVVVVURERFVVVURERERERERERERERERERERERERERDMzMzMzMzMzM1VVVVVVVVVVVURERERERERERERERDMzM0RERDMzM0RERERERDMzM0RERERERERERERERDMzM0RERERERERERFVVVVVVVVVVVURERERERERERERERERERERERERERERERERERERERDMzM0RERCIiIjMzMzMzM0RERERERERERFVVVURERERERERERDMzM0RERDMzM0RERDMzM0RERERERERERERERERERERERERERDMzMzMzMzMzMzMzM0RERFVVVVVVVURERERERDMzMzMzMzMzMzMzMzMzM0RERDMzM0RERDMzMzMzM0RERDMzMzMzMzMzMyIiIiIiIiIiIjMzM0RERFVVVVVVVURERDMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERDMzM0RERHd3d4iIiHd3d0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIkRERERERERERERERERERERERFVVVURERERERERERERERERERERERERERFVVVVVVVURERERERERERERERERERERERFVVVVVVVVVVVWZmZlVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVURERFVVVURERERERFVVVVVVVVVVVURERERERERERERERERERERERERERERERERERERERERERERERERERFVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVURERFVVVWZmZnd3d3d3d3d3d3d3d2ZmZnd3d3d3d2ZmZnd3d3d3d3d3d4iIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZmZmZnd3d3d3d4iIiHd3d3d3d4iIiHd3d3d3d4iIiIiIiJmZmYiIiIiIiIiIiIiIiIiIiJmZmYiIiHd3d2ZmZmZmZmZmZmZmZlVVVURERFVVVVVVVWZmZlVVVWZmZmZmZmZmZlVVVURERDMzMzMzM0RERDMzMzMzMzMzMyIiIjMzMzMzM0RERIiIiMzMzMzMzLu7u6qqqqqqqpmZmZmZmYiIiGZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVURERERERERERERERERERERERDMzM0RERERERERERERERERERERERDMzM0RERERERERERDMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM0RERDMzM0RERERERDMzM0RERCIiIjMzM0RERERERFVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVWZmZlVVVVVVVTMzMzMzMzMzMzMzM0RERGZmZlVVVVVVVURERFVVVWZmZlVVVURERFVVVXd3d2ZmZmZmZlVVVVVVVWZmZnd3d2ZmZlVVVVVVVURERERERERERERERERERGZmZnd3d3d3d0RERERERERERDMzMzMzM0RERERERERERERERERERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERDMzM0RERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVWZmZlVVVVVVVWZmZlVVVVVVVVVVVWZmZnd3d3d3d4iIiIiIiIiIiIiIiJmZmYiIiIiIiIiIiHd3d3d3d3d3d4iIiIiIiJmZmYiIiIiIiGZmZnd3d2ZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiJmZmaqqqpmZmZmZmZmZmYiIiGZmZmZmZlVVVVVVVWZmZnd3d4iIiJmZmczMzN3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////u7u7u7u7u7u7u7u7d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7////u7u7u7u7u7u7d3d3d3d3d3d3MzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7u7u7vMzMzMzMzd3d3MzMzMzMzMzMy7u7vMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7uqqqqqqqqZmZmqqqqZmZmZmZl3d3d3d3d3d3dVVVVERERVVVVERERERERERERERERERERERERERERERERERERERERERERVVVVVVVVERERVVVVERERmZmZmZmZmZmZVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVERERVVVVmZmZ3d3dVVVVmZmZ3d3eIiIhmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVEREQzMzNERERERERERERERERVVVVmZmZVVVVERERVVVVERERERERERERVVVVmZmZVVVVmZmZERERVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERmZmaIiIhmZmZVVVVmZmaIiIh3d3d3d3eZmZmZmZl3d3dmZmZVVVVVVVVmZmZmZmZ3d3dmZmZmZmZ3d3dmZmZVVVVVVVVVVVVVVVVmZmZ3d3dVVVVERERERERmZmZmZmZ3d3eIiIhmZmZVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVERERVVVVmZmZmZmZmZmZmZmZ3d3eIiIi7u7u7u7vd3d3d3d3d3d3u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzd3d3MzMy7u7vd3d3d3d3d3d3MzMzMzMy7u7uqqqqqqqqqqqqqqqqqqqqZmZmZmZl3d3dmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZmZmZ3d3d3d3dmZmZmZmZmZmZmZmZmZmZ3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVV3d3d3d3dmZmZmZmZVVVVVVVVmZmZVVVVVVVVERERVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3dVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZVVVVmZmZVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZ3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVV3d3dmZmZVVVVERERVVVVVVVVVVVVEREREREQzMzMzMzMzMzMzMzNEREREREQzMzNERERERERmZmZ3d3dmZmZmZmZVVVVERERERERVVVVERERERERVVVVVVVVERERVVVVEREREREREREREREREREQzMzNERERmZmZVVVVERERVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVERERVVVVEREREREREREREREQzMzNEREQzMzNVVVVVVVVVVVVEREREREREREREREREREREREREREQzMzMzMzNEREREREQzMzNERERERERERERVVVUzMzNERERERERVVVVVVVVVVVVERERERERERERERERERERERERVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzNERERVVVVVVVVEREREREREREREREREREQzMzNEREREREREREQzMzNEREREREREREREREREREREREQzMzMzMzMzMzNERERVVVVVVVVEREQzMzMzMzNEREQzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIREREiIiIzMzNERERVVVVERERERERERERVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzMiIiIzMzMzMzMiIiIzMzMzMzNEREQzMzMzMzNERESIiIiIiIhVVVUiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzNEREQzMzNEREREREQzMzNEREQzMzNEREREREQzMzNERERERERERERERERERERERERERERERERERERERERERERERERERERVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERVVVVERERERERVVVVERERVVVVVVVVVVVVERERERERERERERERERERVVVVVVVVVVVVmZmZ3d3dmZmZmZmZVVVVmZmZVVVVVVVVVVVVmZmZ3d3eIiIh3d3dmZmZmZmZ3d3dmZmZmZmZmZmZVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3eIiIh3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIh3d3d3d3d3d3eIiIiIiIiIiIiZmZmZmZmIiIh3d3dVVVVmZmZmZmZmZmZVVVVERERVVVVVVVVERERERERERERmZmZVVVVEREQzMzMzMzNVVVVEREQzMzMiIiIzMzMiIiIzMzMzMzNERER3d3e7u7vd3d27u7u7u7uqqqqZmZmZmZl3d3dmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVV3d3dmZmZERERERERERERERERVVVVEREREREREREQzMzNEREREREREREQzMzNEREQzMzMzMzNERERVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNERERERERVVVVEREQzMzMzMzNERERVVVVVVVVVVVVVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVERERERERERERERERVVVVmZmZmZmZVVVVVVVVERERERERmZmZVVVVERERVVVVVVVVmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVEREREREREREREREREREQzMzNERERVVVVVVVVEREREREREREREREQzMzNERERERERERERERERERERERERERERVVVVERERVVVVVVVVVVVVmZmZVVVVVVVVERERVVVVERERERERVVVVERERERERERERVVVVERERVVVVERERVVVVVVVVVVVVVVVVERERVVVVmZmZ3d3dmZmZVVVVVVVVVVVVVVVVVVVVmZmaIiIiZmZmIiIiIiIiIiIh3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIh3d3d3d3eIiIh3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiZmZmZmZmqqqqqqqqqqqqqqqqqqqqZmZmZmZl3d3d3d3d3d3dmZmaIiIiZmZmqqqq7u7vd3d3u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u////7u7u////7u7u7u7u3d3d3d3d3d3dzMzMzMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7zMzMzMzM3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7zMzMzMzMu7u7u7u7qqqqqqqqqqqqmZmZmZmZiIiIiIiId3d3d3d3ZmZmVVVVREREVVVVREREREREREREREREREREREREREREREREREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmVVVVVVVVZmZmd3d3d3d3VVVVZmZmZmZmd3d3d3d3ZmZmZmZmd3d3ZmZmZmZmVVVVREREREREREREVVVVREREMzMzREREREREREREREREREREVVVVVVVVZmZmVVVVVVVVZmZmVVVVREREREREVVVVVVVVVVVVZmZmd3d3d3d3ZmZmVVVVVVVVZmZmVVVVVVVVVVVVVVVVZmZmVVVVREREMzMzREREVVVVVVVVVVVVREREVVVVZmZmd3d3ZmZmVVVVZmZmd3d3d3d3d3d3iIiId3d3d3d3d3d3ZmZmZmZmd3d3ZmZmZmZmVVVVd3d3iIiId3d3VVVVREREREREZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmiIiId3d3ZmZmVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmVVVVZmZmVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmd3d3iIiIqqqqzMzM3d3d7u7u7u7u////7u7u////7u7u7u7u7u7u7u7u3d3d3d3dzMzM3d3dzMzMzMzMzMzM3d3d3d3dzMzMzMzMzMzMu7u7u7u7u7u7mZmZmZmZiIiIiIiIiIiId3d3d3d3ZmZmVVVVREREMzMzREREREREREREREREREREREREREREVVVVREREVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVZmZmd3d3ZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmVVVVVVVVZmZmVVVVZmZmVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmd3d3d3d3d3d3d3d3ZmZmd3d3d3d3ZmZmZmZmZmZmZmZmVVVVVVVVZmZmVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmd3d3d3d3ZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVREREVVVVREREREREREREVVVVREREREREVVVVREREZmZmd3d3iIiId3d3ZmZmVVVVVVVVVVVVVVVVREREREREREREREREREREREREREREREREREREVVVVd3d3mZmZd3d3d3d3REREMzMzREREREREREREREREREREVVVVVVVVREREREREREREREREREREMzMzMzMzREREVVVVZmZmVVVVVVVVVVVVREREVVVVVVVVREREVVVVVVVVVVVVREREVVVVREREREREREREREREREREMzMzREREVVVVVVVVREREREREMzMzREREMzMzREREMzMzREREREREREREREREREREREREREREREREVVVVMzMzREREREREREREVVVVVVVVREREREREVVVVVVVVVVVVVVVVREREVVVVVVVVREREREREMzMzMzMzREREMzMzREREVVVVVVVVREREREREREREREREREREREREREREMzMzREREREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzREREVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzREREREREVVVVREREREREREREREREMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzREREREREMzMzMzMzIiIiREREREREREREIiIiMzMzMzMzMzMzZmZmiIiId3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREREREVVVVVVVVZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVREREREREREREREREREREREREVVVVREREREREVVVVVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmVVVVREREREREVVVVVVVViIiImZmZmZmZiIiId3d3iIiIiIiImZmZiIiId3d3VVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3iIiId3d3d3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3ZmZmZmZmZmZmd3d3ZmZmZmZmd3d3ZmZmd3d3d3d3iIiIiIiIiIiId3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVd3d3d3d3d3d3iIiIiIiIiIiId3d3iIiIiIiIiIiImZmZmZmZiIiIiIiId3d3ZmZmZmZmZmZmZmZmZmZmREREVVVVZmZmREREREREMzMzREREZmZmVVVVMzMzMzMzMzMzVVVVREREMzMzIiIiMzMzMzMzMzMzMzMzREREZmZmu7u7zMzMzMzMqqqqmZmZd3d3mZmZd3d3ZmZmVVVVZmZmd3d3ZmZmVVVVVVVVd3d3ZmZmZmZmVVVVREREREREVVVVVVVVREREMzMzREREMzMzMzMzREREREREMzMzMzMzMzMzVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREVVVVVVVVVVVVREREREREREREREREVVVVVVVVVVVVREREREREREREREREVVVVREREVVVVREREREREREREVVVVd3d3iIiId3d3VVVVVVVVREREREREVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVREREREREVVVVREREREREREREMzMzMzMzMzMzREREMzMzMzMzREREMzMzMzMzREREREREREREREREMzMzREREREREREREREREVVVVREREREREREREVVVVd3d3d3d3ZmZmVVVVREREREREREREREREREREVVVVREREVVVVREREREREVVVVREREVVVVREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmd3d3d3d3iIiId3d3ZmZmZmZmd3d3ZmZmd3d3d3d3d3d3d3d3ZmZmiIiId3d3iIiIiIiImZmZmZmZiIiIiIiImZmZmZmZiIiId3d3d3d3iIiId3d3d3d3d3d3iIiIiIiIiIiImZmZiIiIiIiImZmZmZmZqqqqmZmZqqqqqqqqqqqqqqqqqqqqiIiIiIiImZmZmZmZmZmZqqqqzMzMzMzM3d3d////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7v///+7u7u7u7u7u7t3d3d3d3e7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3czMzMzMzMzMzLu7u8zMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u8zMzN3d3d3d3d3d3czMzMzMzN3d3czMzN3d3czMzN3d3czMzLu7u7u7u7u7u7u7u6qqqqqqqqqqqqqqqpmZmZmZmZmZmXd3d3d3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVURERERERERERERERERERFVVVVVVVVVVVWZmZlVVVVVVVURERFVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d3d3d2ZmZlVVVVVVVVVVVVVVVVVVVWZmZnd3d2ZmZmZmZmZmZnd3d3d3d3d3d2ZmZnd3d2ZmZlVVVVVVVURERERERCIiIjMzMzMzMzMzM0RERFVVVVVVVVVVVWZmZmZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVURERERERERERERERERERERERFVVVVVVVWZmZnd3d1VVVVVVVWZmZmZmZnd3d2ZmZlVVVWZmZmZmZmZmZnd3d2ZmZmZmZmZmZnd3d3d3d3d3d1VVVVVVVVVVVXd3d3d3d3d3d2ZmZkRERERERFVVVVVVVVVVVVVVVXd3d3d3d2ZmZmZmZnd3d2ZmZmZmZkRERFVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZnd3d5mZmczMzN3d3e7u7v///////////+7u7v///////+7u7v///+7u7u7u7u7u7t3d3d3d3czMzLu7u7u7u8zMzN3d3d3d3d3d3bu7u5mZmaqqqqqqqpmZmYiIiHd3d3d3d2ZmZmZmZmZmZlVVVURERDMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERDMzM0RERDMzM0RERERERERERFVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVVVVVWZmZmZmZnd3d2ZmZmZmZmZmZlVVVVVVVURERGZmZlVVVVVVVWZmZmZmZnd3d2ZmZmZmZkRERERERFVVVWZmZmZmZlVVVWZmZlVVVWZmZlVVVWZmZmZmZmZmZlVVVWZmZmZmZnd3d3d3d2ZmZmZmZnd3d3d3d2ZmZmZmZlVVVURERFVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVURERFVVVWZmZlVVVWZmZmZmZnd3d3d3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVXd3d3d3d4iIiIiIiHd3d1VVVVVVVWZmZlVVVURERFVVVVVVVVVVVVVVVVVVVVVVVURERERERGZmZpmZmZmZmYiIiHd3d1VVVURERDMzM0RERERERFVVVURERERERERERFVVVURERERERERERERERDMzM0RERERERFVVVWZmZlVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVURERERERERERERERFVVVURERERERDMzM0RERERERFVVVVVVVVVVVURERERERERERDMzM0RERERERDMzM0RERERERERERERERFVVVURERFVVVURERDMzM0RERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERDMzMzMzMzMzM0RERERERFVVVVVVVURERERERERERERERDMzM0RERERERERERERERERERDMzM0RERDMzM0RERERERDMzMyIiIjMzMyIiIjMzM0RERFVVVURERERERDMzMzMzM0RERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzM0RERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERDMzMzMzMzMzM2ZmZmZmZjMzMyIiIjMzMzMzMzMzM2ZmZoiIiGZmZkRERERERERERERERDMzMzMzMzMzM0RERERERFVVVWZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERERERERERERERERERFVVVURERERERFVVVVVVVVVVVVVVVURERFVVVURERERERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZlVVVWZmZnd3d2ZmZnd3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVURERFVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERFVVVYiIiJmZmZmZmZmZmYiIiIiIiIiIiJmZmYiIiHd3d2ZmZlVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d3d3d3d3d3d3d4iIiHd3d2ZmZmZmZnd3d3d3d3d3d3d3d2ZmZnd3d2ZmZnd3d2ZmZnd3d4iIiIiIiIiIiJmZmYiIiIiIiIiIiIiIiJmZmZmZmYiIiHd3d3d3d2ZmZmZmZmZmZnd3d1VVVURERGZmZmZmZkRERDMzM0RERFVVVWZmZlVVVTMzMyIiIjMzM0RERERERCIiIjMzMzMzMyIiIjMzMzMzM0RERFVVVaqqqt3d3bu7u6qqqoiIiIiIiIiIiIiIiGZmZlVVVVVVVWZmZmZmZlVVVWZmZoiIiGZmZlVVVVVVVURERFVVVVVVVVVVVURERERERDMzM0RERFVVVURERDMzMzMzMzMzM0RERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERERERFVVVVVVVURERERERERERERERFVVVWZmZlVVVURERFVVVVVVVURERERERERERERERERERERERFVVVWZmZpmZmYiIiGZmZkRERERERERERFVVVURERERERFVVVVVVVURERERERERERFVVVVVVVVVVVVVVVURERERERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERERERERERERERERERFVVVURERERERFVVVWZmZnd3d3d3d2ZmZkRERERERERERERERERERERERERERFVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVVVVVURERFVVVWZmZmZmZlVVVVVVVXd3d3d3d2ZmZlVVVWZmZmZmZmZmZnd3d3d3d4iIiHd3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiJmZmZmZmZmZmZmZmZmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d4iIiIiIiJmZmaqqqqqqqqqqqqqqqqqqqqqqqoiIiIiIiJmZmaqqqqqqqszMzMzMzO7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3u7u7d3d3u7u7d3d3d3d3d3d3MzMy7u7u7u7u7u7vMzMzMzMzMzMzMzMzd3d3MzMzMzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7uqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqZmZl3d3d3d3dmZmZVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZmZmZVVVVVVVVERERVVVVVVVVERERVVVVVVVVmZmZmZmZ3d3dmZmZmZmZVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVEREQzMzNEREQzMzMzMzMzMzMzMzNERERVVVVVVVVmZmZmZmZVVVVVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZ3d3dmZmZmZmZVVVVVVVVERERVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZmZmZ3d3d3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3dVVVVVVVVmZmZ3d3dmZmZmZmZ3d3d3d3dVVVUzMzNVVVV3d3dVVVVmZmZ3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERVVVVmZmZ3d3dmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZ3d3eqqqq7u7vd3d3////u7u7////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3MzMyZmZmIiIiqqqrMzMy7u7uZmZlmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZ3d3dmZmZmZmZVVVVEREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERVVVVVVVVVVVVmZmZmZmZ3d3eIiIh3d3eIiIh3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZ3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVERERERERVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZVVVVmZmZmZmZVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVmZmZVVVVVVVVVVVVVVVVmZmZ3d3eIiIiIiIiIiIh3d3dmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3eIiIiqqqqZmZmIiIh3d3dVVVVERERERERERERVVVVERERVVVVVVVVVVVVVVVVVVVVEREREREREREREREQzMzNERERVVVVmZmZVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVERERVVVVEREREREREREREREQzMzMzMzNVVVVmZmZVVVVEREQzMzNEREREREQzMzNERERERERVVVVERERVVVVERERVVVVERERVVVVEREREREQzMzNVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZVVVVVVVVmZmZVVVVVVVVVVVVEREREREREREQzMzNERERVVVVVVVVVVVVERERERERERERERERVVVVVVVVVVVVEREREREREREQzMzNEREQzMzNEREREREQzMzMiIiIzMzMiIiJERERVVVVVVVVEREREREQzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMiIiIiIiIREREiIiIzMzNEREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNmZmaIiIhVVVUiIiIzMzMzMzNEREQzMzNERER3d3eIiIhmZmZVVVVVVVVVVVVVVVVERERERERVVVVVVVVmZmZmZmZVVVVVVVVVVVVERERERERVVVVERERVVVVERERVVVVERERVVVVEREREREREREREREREREREREREREREREQzMzNEREQzMzNERERVVVVERERERERERERVVVVERERVVVVERERVVVVERERERERERERVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZVVVVmZmZVVVVmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3dmZmZ3d3dmZmZ3d3dmZmZ3d3d3d3d3d3dmZmZ3d3dmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3dmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3dmZmZmZmZmZmZVVVVVVVVmZmZVVVVVVVVERERVVVVERERVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZ3d3dmAP//AABmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZnd3d3d3d4iIiHd3d3d3d3d3d3d3d3d3d2ZmZnd3d4iIiJmZmZmZmYiIiIiIiJmZmaqqqpmZmZmZmXd3d2ZmZlVVVWZmZoiIiGZmZkRERERERGZmZlVVVURERDMzM0RERHd3d2ZmZkRERDMzMzMzMzMzM0RERERERDMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERJmZmczMzLu7u6qqqoiIiIiIiIiIiIiIiFVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d2ZmZlVVVVVVVURERFVVVURERFVVVURERERERDMzMzMzM1VVVVVVVURERDMzMzMzMzMzM0RERFVVVURERERERDMzM0RERERERERERERERERERDMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERFVVVURERERERERERERERFVVVURERFVVVVVVVVVVVURERFVVVURERFVVVURERERERFVVVVVVVVVVVZmZmaqqqnd3d1VVVURERERERDMzM0RERERERERERERERFVVVURERERERERERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERERERDMzM0RERFVVVURERERERERERFVVVURERDMzM0RERERERERERERERERERERERERERFVVVVVVVVVVVURERFVVVURERERERERERERERERERFVVVURERERERFVVVURERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d2ZmZnd3d2ZmZmZmZmZmZnd3d3d3d4iIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d4iIiJmZmZmZmZmZmZmZmZmZmYiIiJmZmZmZmZmZmZmZmYiIiHd3d3d3d3d3d2ZmZnd3d3d3d4iIiIiIiKqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqru7u8zMzN3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3MzMzMzMzMzMzMzMzMzMzd3d3u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3MzMzMzMzMzMy7u7vMzMy7u7vMzMzMzMy7u7vMzMy7u7vMzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7uqqqq7u7uqqqq7u7uqqqqqqqqZmZmZmZmZmZmIiIiIiIiIiIh3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVV3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3dmZmZmZmZmZmZVVVVVVVVEREQzMzMzMzNEREREREREREQzMzNERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZ3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVmZmZmZmZmZmZmZmZ3d3eIiIh3d3d3d3d3d3d3d3eIiIiIiIiZmZmIiIh3d3d3d3d3d3d3d3dVVVVVVVV3d3d3d3dmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZVVVVVVVVVVVVmZmZVVVVERERVVVVVVVVERERERERVVVVmZmZ3d3dmZmZVVVVVVVVmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZ3d3eqqqrMzMzu7u7u7u7////u7u7u7u7u7u7u7u7u7u7d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7MzMy7u7uZmZmIiIiqqqqqqqqqqqpmZmZVVVVmZmZERERVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZ3d3d3d3d3d3dmZmZ3d3dVVVVVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzNERERERERERERVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZVVVVVVVVmZmZmZmZVVVVVVVVERERERERVVVVVVVVERERVVVVVVVVmZmZmZmZVVVVmZmZmZmZmZmZVVVVmZmZVVVVVVVVmZmZmZmZVVVVVVVVVVVVmZmZVVVVVVVVERERVVVVERERVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZ3d3dmZmZmZmZmZmZ3d3d3d3d3d3d3d3dVVVVERERVVVVERERVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3d3d3d3d3eIiIh3d3dmZmZ3d3dmZmZ3d3d3d3d3d3dmZmZ3d3d3d3d3d3eIiIiIiIiZmZmZmZmIiIiZmZmZmZmqqqqZmZl3d3dEREQzMzNERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERERERVVVVmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVEREREREQzMzMzMzNERERVVVVmZmZVVVVEREREREREREQzMzNERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVmZmZ3d3dmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZ3d3d3d3dmZmZVVVVEREREREQzMzNERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVEREREREREREREREREREQzMzMzMzMzMzMzMzMzMzNERERVVVVVVVVEREQzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMiIiIiIiIiIiIzMzMiIiIzMzMzMzNEREREREREREQzMzNEREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiJEREREREQzMzMzMzMzMzNEREQzMzMzMzMzMzNERERmZmZmZmYzMzNERERERERVVVVERERERERERERERERERERERERERERERERERERVVVVERERVVVVVVVVEREREREREREREREREREREREREREREREQzMzNERERERERERERERERERERERERERERERERERERVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZVVVVmZmZVVVVmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZmZmZ3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIh3d3d3d3d3d3eIiIiIiIh3d3eIiIh3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIiZmZl3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZ3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZVVVVmZmZVVVVmZmZVVVVVVVVmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3eIiIiIiIiZmZmZmZmZmZmZmZmZmZmZmZmZmZmqqqqZmZlVVVVVVVVVVVVmZmZ3d3dVVVVERERmZmZmZmZEREREREQzMzNVVVWIiIhmZmZEREQzMzMzMzMiIiIzMzNEREQzMzMiIiIzMzMzMzMiIiIzMzMzMzNVVVWZmZnMzMzMzMyqqqqIiIiIiIiIiIh3d3dmZmZERERVVVVVVVVVVVVmZmaIiIhmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVERERERERVVVVERERERERVVVVVVVVEREQzMzNERERERERVVVVVVVVEREREREREREREREREREREREREREQzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzNERERERERERERVVVVVVVVERERERERERERERERERERERERVVVVVVVVERERVVVVVVVVmZmZmZmaIiIiZmZmIiIhmZmZVVVVEREQzMzMzMzNEREREREQzMzNERERERERVVVVVVVVVVVVERERVVVVVVVVmZmZ3d3d3d3dVVVVVVVVmZmZERERERERERERERERVVVVVVVVERERERERERERERERERERERERERERERERERERVVVVERERVVVVVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVEREREREREREQzMzNVVVVERERVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmZ3d3dmZmZ3d3d3d3eIiIiZmZmIiIh3d3d3d3eIiIh3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3eIiIiIiIiZmZmZmZmZmZmZmZmZmZmIiIiIiIh3d3d3d3dmZmZmZmZVVVVVVVVmZmZ3d3d3d3eIiIiZmZmZmZmZmZmqqqqqqqq7u7u7u7vMzMzMzMzd3d3d3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u7u7u////7u7u7u7u////7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3dzMzM3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzMu7u7u7u7u7u7u7u7u7u7qqqqqqqqu7u7zMzMu7u7zMzMzMzMzMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7qqqqu7u7qqqqmZmZu7u7qqqqmZmZmZmZd3d3d3d3d3d3ZmZmd3d3d3d3VVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVREREVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVREREREREMzMzREREREREREREREREVVVVREREREREREREREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmd3d3ZmZmZmZmd3d3ZmZmVVVVREREREREVVVVVVVVVVVVVVVVZmZmVVVVZmZmREREVVVVVVVVVVVVVVVVVVVVZmZmd3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiId3d3iIiId3d3d3d3d3d3iIiId3d3d3d3ZmZmZmZmZmZmd3d3VVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVREREREREVVVVREREVVVVZmZmVVVVVVVVVVVVZmZmVVVVVVVVVVVVZmZmZmZmVVVVVVVVREREZmZmiIiImZmZmZmZzMzM3d3d////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u7u7uzMzMu7u7u7u7qqqqu7u7qqqqiIiId3d3iIiId3d3d3d3ZmZmZmZmiIiIZmZmZmZmVVVVZmZmZmZmd3d3VVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVREREREREREREMzMzMzMzMzMzMzMzREREMzMzREREMzMzREREREREREREREREVVVVZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiId3d3d3d3ZmZmZmZmd3d3ZmZmREREREREVVVVREREVVVVREREREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVREREVVVVVVVVZmZmZmZmVVVVREREVVVVREREVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmd3d3ZmZmVVVVREREREREVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVZmZmd3d3d3d3d3d3d3d3d3d3iIiId3d3ZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiImZmZmZmZmZmZqqqqqqqqqqqqmZmZd3d3VVVVREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmVVVVREREREREVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3ZmZmZmZmZmZmVVVVVVVVREREREREREREMzMzREREVVVVVVVVREREREREREREREREREREREREVVVVZmZmVVVVZmZmVVVVZmZmVVVVZmZmVVVVVVVVVVVVREREZmZmd3d3ZmZmZmZmd3d3d3d3ZmZmd3d3d3d3ZmZmZmZmd3d3d3d3ZmZmVVVVREREREREMzMzMzMzVVVVVVVVVVVVREREREREVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVREREREREREREREREREREMzMzMzMzIiIiMzMzMzMzVVVVREREREREMzMzREREREREREREMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiREREREREREREREREMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzIiIiMzMzMzMzIiIiIiIiMzMzMzMzMzMzREREMzMzMzMzMzMzVVVVREREREREMzMzREREMzMzREREMzMzREREMzMzREREREREREREREREREREREREREREREREVVVVVVVVVVVVREREVVVVREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmd3d3d3d3ZmZmd3d3ZmZmd3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3iIiId3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZmZmZiIiIiIiIiIiIiIiId3d3iIiId3d3iIiId3d3iIiIiIiId3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiId3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3iIiIiIiId3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmd3d3iIiImZmZmZmZqqqqqqqqqqqqmZmZmZmZiIiIqqqqmZmZiIiIZmZmREREREREd3d3d3d3REREREREd3d3ZmZmMzMzMzMzREREREREZmZmVVVVREREREREMzMzIiIiMzMzREREMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREiIiIzMzMzMzMqqqqmZmZiIiId3d3iIiIZmZmVVVVREREVVVVZmZmd3d3d3d3VVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVREREREREREREREREVVVVVVVVREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREMzMzREREREREMzMzMzMzVVVVREREREREREREREREVVVVREREREREREREREREREREREREREREVVVVREREVVVVVVVVZmZmiIiImZmZiIiId3d3VVVVMzMzREREMzMzMzMzMzMzREREMzMzMzMzREREREREZmZmZmZmVVVVVVVVVVVVVVVVd3d3d3d3ZmZmVVVVVVVVVVVVREREVVVVREREVVVVVVVVVVVVMzMzREREREREVVVVVVVVREREREREVVVVZmZmVVVVVVVVVVVVREREVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVREREREREREREVVVVREREREREVVVVREREREREVVVVVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmZmZmd3d3ZmZmd3d3d3d3iIiIiIiIiIiId3d3d3d3iIiId3d3ZmZmVVVVZmZmVVVVVVVVZmZmZmZmd3d3d3d3iIiImZmZmZmZqqqqmZmZmZmZiIiId3d3ZmZmZmZmVVVVVVVVZmZmZmZmZmZmZmZmd3d3iIiIiIiImZmZmZmZqqqqqqqqu7u7u7u7zMzM3d3d3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7u7u7u7u7t3d3e7u7u7u7u7u7u7u7t3d3d3d3d3d3czMzMzMzLu7u7u7u7u7u6qqqru7u7u7u7u7u7u7u8zMzMzMzMzMzLu7u8zMzMzMzLu7u8zMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u6qqqru7u6qqqqqqqqqqqpmZmYiIiIiIiHd3d3d3d2ZmZmZmZkRERERERERERERERFVVVURERFVVVVVVVWZmZmZmZnd3d3d3d2ZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZlVVVVVVVURERERERERERERERERERFVVVVVVVVVVVURERFVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d4iIiHd3d2ZmZmZmZmZmZmZmZlVVVVVVVURERERERERERERERERERFVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d4iIiJmZmYiIiIiIiIiIiHd3d4iIiHd3d3d3d3d3d3d3d3d3d4iIiJmZmaqqqoiIiGZmZlVVVWZmZmZmZmZmZlVVVVVVVVVVVWZmZlVVVVVVVURERFVVVURERERERERERERERFVVVVVVVWZmZmZmZlVVVVVVVVVVVURERFVVVVVVVVVVVWZmZkRERERERERERGZmZpmZmczMzN3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7v///+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7v///+7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3czMzMzMzLu7u6qqqoiIiGZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVURERFVVVURERERERERERERERERERFVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVURERERERERERERERERERFVVVVVVVVVVVWZmZnd3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d4iIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d2ZmZkRERERERERERERERFVVVURERFVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVXd3d2ZmZlVVVVVVVURERERERERERERERFVVVVVVVWZmZlVVVVVVVVVVVWZmZmZmZmZmZoiIiHd3d1VVVVVVVWZmZmZmZnd3d2ZmZkRERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d4iIiHd3d4iIiIiIiIiIiHd3d2ZmZlVVVWZmZmZmZmZmZmZmZnd3d4iIiHd3d4iIiIiIiIiIiJmZmZmZmZmZmaqqqru7u6qqqoiIiGZmZlVVVURERFVVVVVVVVVVVWZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d2ZmZlVVVURERERERFVVVXd3d2ZmZlVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZnd3d2ZmZmZmZmZmZmZmZlVVVVVVVURERERERERERGZmZlVVVURERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVWZmZlVVVVVVVURERFVVVWZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZnd3d2ZmZnd3d1VVVVVVVURERERERERERERERFVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVURERERERDMzMzMzMzMzMzMzMyIiIkRERERERERERERERDMzM0RERERERERERDMzM0RERDMzM0RERDMzMzMzMzMzM0RERDMzMzMzMyIiIjMzMyIiIjMzMzMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIjMzM0RERERERERERCIiIjMzMzMzM0RERERERERERERERERERERERERERERERERERFVVVURERERERERERERERFVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVURERERERERERFVVVVVVVVVVVVVVVWZmZmZmZlVVVWZmZmZmZnd3d2ZmZnd3d3d3d2ZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZlVVVVVVVWZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZlVVVWZmZlVVVWZmZlVVVWZmZlVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZoiIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiIiIiHd3d4iIiHd3d3d3d3d3d3d3d4iIiHd3d4iIiHd3d3d3d3d3d4iIiIiIiHd3d4iIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZmZmZnd3d2ZmZnd3d3d3d2ZmZnd3d2ZmZnd3d3d3d4iIiIiIiHd3d3d3d2ZmZnd3d2ZmZnd3d3d3d5mZmZmZmaqqqqqqqpmZmZmZmZmZmZmZmZmZmaqqqoiIiHd3d1VVVURERFVVVWZmZlVVVURERFVVVWZmZlVVVTMzM0RERERERERERFVVVWZmZkRERDMzMzMzMzMzMyIiIjMzMzMzMyIiIiIiIjMzMzMzMzMzM0RERERERHd3d7u7u7u7u6qqqpmZmYiIiIiIiHd3d3d3d2ZmZlVVVVVVVWZmZnd3d1VVVURERFVVVVVVVWZmZlVVVVVVVVVVVVVVVURERERERFVVVVVVVURERFVVVVVVVWZmZlVVVURERFVVVVVVVVVVVWZmZmZmZmZmZlVVVURERERERERERERERERERDMzM0RERDMzM0RERERERFVVVURERERERERERERERERERDMzM0RERERERERERERERFVVVURERFVVVVVVVVVVVVVVVXd3d4iIiIiIiHd3d1VVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERFVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVVVVVURERERERERERERERERERFVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVURERFVVVURERFVVVXd3d2ZmZmZmZnd3d2ZmZlVVVWZmZnd3d4iIiHd3d2ZmZmZmZnd3d3d3d2ZmZnd3d3d3d3d3d3d3d4iIiHd3d2ZmZmZmZmZmZlVVVWZmZmZmZoiIiIiIiJmZmZmZmZmZmZmZmZmZmYiIiHd3d2ZmZlVVVVVVVVVVVWZmZmZmZnd3d3d3d3d3d4iIiIiIiJmZmZmZmaqqqru7u7u7u8zMzN3d3e7u7u7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3MzMzMzMy7u7u7u7u7u7u7u7vMzMy7u7uqqqq7u7uqqqq7u7u7u7vMzMy7u7vMzMzMzMzMzMzMzMzd3d3MzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7uqqqq7u7uqqqqqqqqqqqqZmZmZmZmIiIhmZmZmZmZVVVVVVVVERERERERERERVVVVVVVVVVVVmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3dmZmZ3d3d3d3dmZmZmZmZmZmZVVVVERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZ3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3eIiIiIiIh3d3d3d3dmZmZVVVVVVVVVVVVEREREREREREQzMzMzMzNVVVVERERERERVVVVVVVVVVVVVVVVmZmZmZmZVVVV3d3d3d3eIiIiIiIh3d3eIiIiZmZmZmZmIiIiIiIh3d3d3d3dmZmZmZmZmZmZ3d3d3d3d3d3eIiIiZmZmZmZmIiIhmZmZVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZEREREREREREREREREREQzMzNERERVVVVmZmZVVVVmZmZVVVVVVVVVVVVERERVVVVVVVVERERERERERERERERmZmaZmZnMzMzu7u7////////////////u7u7u7u7u7u7////u7u7u7u7////u7u7u7u7////u7u7u7u7u7u7u7u7u7u7MzMzd3d3MzMy7u7u7u7u7u7u7u7u7u7uqqqqqqqqZmZmIiIhmZmZERERERERVVVVEREREREREREREREREREREREQzMzNEREQzMzNEREREREREREREREREREREREREREREREQzMzNEREQzMzNERERERERVVVVmZmZmZmZ3d3eIiIh3d3d3d3d3d3dmZmZVVVVERERVVVVVVVVERERVVVVVVVV3d3eIiIh3d3d3d3eIiIiZmZmIiIh3d3dmZmZmZmZmZmZmZmZmZmaIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIiIiIh3d3dmZmZVVVVERERERERERERERERERERVVVVVVVVmZmZmZmZ3d3dmZmZmZmZ3d3d3d3dmZmZmZmZmZmZmZmZVVVVVVVVmZmZ3d3dVVVVVVVVVVVVERERERERERERERERERERVVVVVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZVVVVmZmZmZmZ3d3d3d3dmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3dmZmZ3d3eZmZmZmZmIiIh3d3eIiIh3d3dVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3eIiIiZmZmIiIiIiIiZmZmqqqqqqqq7u7uqqqp3d3dVVVVERERERERVVVVVVVVVVVVmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3dmZmZmZmZVVVVERERVVVVmZmZmZmZVVVVERERERERVVVVmZmZVVVVmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3dmZmZVVVVERERERERERERVVVVmZmZERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVmZmZ3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZ3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZVVVVVVVVmZmZVVVVVVVVEREREREREREQiIiIzMzMiIiIzMzNVVVVERERVVVVEREQzMzNEREREREREREREREREREREREQzMzNEREQzMzMzMzMzMzMzMzMiIiIiIiIzMzMzMzMzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMiIiIzMzMzMzMiIiIiIiIiIiIzMzNEREREREREREQzMzMiIiIzMzNEREREREQzMzMzMzMzMzMzMzMzMzNERERERERERERVVVVERERERERVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVERERERERVVVVERERVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZ3d3d3d3dmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZmZmZmZmZVVVVmZmZVVVVVVVVmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmaIiIiZmZmZmZmZmZmZmZmIiIiIiIiZmZmIiIh3d3eIiIiIiIiIiIiIiIiIiIh3d3dmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3d3d3eIiIh3d3d3d3d3d3d3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZ3d3eIiIiIiIh3d3eIiIh3d3dmZmZmZmZ3d3d3d3eIiIiZmZmZmZmqqqqZmZmqqqqZmZmqqqqZmZmqqqqZmZl3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERERERVVVVERERERERERERVVVVmZmZVVVVERERVVVUzMzMiIiIzMzNEREQzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzNERESqqqrMzMy7u7uqqqqZmZmIiIiIiIiIiIh3d3dVVVVVVVV3d3dVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVEREQzMzMzMzMzMzMzMzNEREQzMzNERERERERVVVVVVVVEREREREREREREREQzMzNEREQzMzNERERERERERERERERERERERERVVVVmZmZmZmZ3d3eIiIhmZmZmZmZEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERVVVVmZmZVVVVmZmZ3d3dmZmZmZmZVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERERERERERERERVVVVERERVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVmZmZmZmZ3d3dVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZ3d3d3d3dmZmZ3d3d3d3dmZmaIiIiIiIh3d3dmZmZVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3eIiIiIiIh3d3d3d3d3d3d3d3eIiIiZmZmqqqqZmZmqqqqqqqqqqqqZmZmIiIh3d3d3d3dmZmZmZmZ3d3d3d3d3d3d3d3eIiIiIiIiZmZmZmZmZmZmqqqq7u7vMzMzd3d3u7u7u7u7u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u7u7u3d3d3d3d3d3d7u7u3d3d3d3d7u7u3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3du7u7u7u7u7u7qqqqmZmZiIiImZmZmZmZqqqqqqqqqqqqu7u7qqqqu7u7u7u7zMzMzMzMzMzMzMzMzMzM3d3dzMzM3d3d3d3dzMzMzMzMu7u7u7u7qqqqqqqqqqqqu7u7u7u7u7u7u7u7u7u7qqqqqqqqmZmZiIiId3d3d3d3VVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVd3d3ZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmVVVVREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3ZmZmd3d3iIiId3d3iIiIiIiId3d3d3d3ZmZmVVVVVVVVREREREREREREREREREREREREREREREREVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVZmZmiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3ZmZmd3d3mZmZiIiIZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVREREREREREREREREREREREREVVVVVVVVZmZmVVVVVVVVREREREREREREVVVVVVVVREREREREVVVVd3d3qqqq3d3d7u7u7u7u////////7u7u////7u7u7u7u7u7u////7u7u////7u7u7u7u////7u7u7u7u7u7u7u7uzMzMqqqqmZmZiIiId3d3d3d3VVVVVVVVZmZmZmZmZmZmVVVVZmZmVVVVREREREREMzMzREREMzMzREREVVVVREREREREVVVVVVVVREREREREMzMzMzMzMzMzMzMzMzMzREREREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREVVVVZmZmd3d3ZmZmd3d3d3d3d3d3d3d3d3d3VVVVZmZmVVVVVVVVVVVVZmZmd3d3iIiIiIiIiIiImZmZmZmZmZmZmZmZiIiIiIiIiIiId3d3iIiIqqqqmZmZiIiId3d3d3d3d3d3iIiId3d3iIiId3d3VVVVREREREREREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVREREREREREREVVVVVVVVREREREREREREVVVVVVVVVVVVZmZmVVVVZmZmVVVVVVVVZmZmZmZmd3d3d3d3d3d3ZmZmVVVVVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVZmZmVVVVVVVVZmZmd3d3ZmZmiIiImZmZd3d3d3d3ZmZmZmZmVVVVVVVVVVVVREREVVVVVVVVZmZmd3d3d3d3iIiId3d3iIiImZmZmZmZmZmZqqqqqqqqqqqqmZmZZmZmVVVVREREREREVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3d3d3iIiId3d3d3d3ZmZmZmZmVVVVVVVVZmZmZmZmZmZmREREREREVVVVVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmd3d3ZmZmZmZmVVVVVVVVZmZmd3d3ZmZmREREREREMzMzREREVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmd3d3d3d3d3d3ZmZmZmZmd3d3d3d3d3d3d3d3d3d3ZmZmZmZmd3d3ZmZmVVVVVVVVVVVVZmZmd3d3iIiIZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVREREREREREREMzMzMzMzIiIiMzMzMzMzREREVVVVVVVVREREREREREREREREMzMzREREMzMzREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzREREREREREREMzMzMzMzMzMzREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREMzMzREREREREREREREREREREREREVVVVREREVVVVVVVVREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmiIiId3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmiIiImZmZqqqqqqqqmZmZmZmZqqqqmZmZmZmZmZmZmZmZiIiIiIiImZmZiIiId3d3ZmZmVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmVVVVZmZmd3d3d3d3ZmZmVVVVZmZmZmZmVVVVZmZmZmZmZmZmd3d3d3d3d3d3ZmZmd3d3ZmZmZmZmZmZmd3d3ZmZmZmZmd3d3ZmZmZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmd3d3iIiImZmZmZmZqqqqqqqqmZmZmZmZqqqqqqqqmZmZd3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVREREREREVVVVVVVVZmZmVVVVREREVVVVVVVVVVVVMzMzREREMzMzMzMzMzMzIiIiMzMzIiIiMzMzREREREREMzMzMzMzREREmZmZzMzMqqqqqqqqqqqqmZmZmZmZmZmZiIiId3d3d3d3d3d3REREREREVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmVVVVMzMzMzMzMzMzMzMzREREREREMzMzMzMzREREVVVVREREREREVVVVVVVVREREMzMzREREREREREREREREREREREREREREMzMzREREVVVVVVVVZmZmd3d3ZmZmREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzREREMzMzREREVVVVVVVVVVVVVVVVZmZmd3d3d3d3d3d3ZmZmVVVVVVVVVVVVVVVVVVVVREREREREVVVVVVVVREREVVVVREREREREREREREREMzMzREREVVVVVVVVd3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3VVVVVVVVZmZmZmZmd3d3d3d3d3d3iIiIiIiIiIiId3d3iIiIiIiId3d3d3d3d3d3ZmZmZmZmVVVVVVVVZmZmVVVVd3d3iIiIiIiIiIiIiIiIiIiId3d3iIiIiIiIiIiImZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZiIiId3d3iIiIiIiIiIiIiIiImZmZmZmZmZmZmZmZmZmZmZmZqqqqu7u7u7u7zMzM3d3d7u7u7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7t3d3bu7u8zMzLu7u8zMzMzMzMzMzN3d3d3d3e7u7t3d3e7u7u7u7u7u7u7u7u7u7szMzLu7u6qqqoiIiHd3d4iIiIiIiIiIiHd3d4iIiJmZmaqqqqqqqqqqqqqqqqqqqqqqqru7u8zMzMzMzMzMzN3d3d3d3czMzMzMzMzMzMzMzLu7u7u7u7u7u6qqqru7u6qqqru7u6qqqru7u6qqqqqqqqqqqqqqqpmZmZmZmYiIiIiIiHd3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d2ZmZmZmZnd3d3d3d2ZmZmZmZnd3d3d3d2ZmZmZmZmZmZlVVVVVVVURERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVWZmZnd3d3d3d2ZmZnd3d3d3d3d3d2ZmZmZmZnd3d3d3d4iIiHd3d3d3d3d3d3d3d4iIiHd3d2ZmZmZmZlVVVVVVVURERERERERERERERFVVVURERFVVVVVVVURERERERERERFVVVURERFVVVVVVVVVVVVVVVWZmZmZmZoiIiJmZmZmZmYiIiIiIiHd3d3d3d2ZmZmZmZnd3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiHd3d2ZmZnd3d4iIiIiIiHd3d2ZmZnd3d3d3d2ZmZlVVVVVVVURERERERERERERERERERERERFVVVVVVVVVVVWZmZlVVVVVVVURERERERFVVVURERFVVVVVVVWZmZnd3d6qqqszMzO7u7v///////////+7u7v///////+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7v///+7u7u7u7szMzJmZmYiIiHd3d2ZmZlVVVVVVVURERFVVVURERFVVVVVVVURERERERDMzM0RERDMzM0RERERERERERERERERERERERFVVVURERFVVVURERERERERERDMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZlVVVWZmZnd3d2ZmZmZmZmZmZnd3d2ZmZnd3d4iIiKqqqqqqqpmZmZmZmXd3d4iIiJmZmaqqqpmZmYiIiHd3d3d3d3d3d3d3d4iIiHd3d2ZmZkRERFVVVURERERERFVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVURERFVVVVVVVVVVVVVVVURERERERERERGZmZlVVVVVVVWZmZlVVVWZmZlVVVWZmZnd3d3d3d3d3d2ZmZmZmZlVVVWZmZlVVVURERERERERERERERFVVVVVVVVVVVVVVVWZmZlVVVWZmZnd3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVURERERERGZmZoiIiIiIiIiIiIiIiJmZmYiIiIiIiIiIiJmZmaqqqpmZmYiIiGZmZkRERERERERERERERERERERERFVVVWZmZnd3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d2ZmZmZmZmZmZmZmZnd3d1VVVVVVVURERFVVVVVVVVVVVVVVVWZmZnd3d3d3d3d3d3d3d3d3d4iIiHd3d1VVVVVVVXd3d3d3d3d3d2ZmZlVVVURERDMzMzMzM0RERERERERERFVVVVVVVVVVVVVVVVVVVXd3d3d3d2ZmZmZmZlVVVWZmZmZmZnd3d2ZmZmZmZlVVVWZmZmZmZnd3d3d3d3d3d3d3d1VVVWZmZmZmZmZmZmZmZmZmZmZmZoiIiJmZmXd3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERERERDMzMzMzMzMzMyIiIiIiIjMzM1VVVURERERERDMzM0RERDMzMzMzM0RERERERERERDMzM0RERDMzM0RERDMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERERERERERDMzM0RERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERDMzMzMzMzMzM0RERERERFVVVURERFVVVURERERERERERERERERERERERFVVVURERFVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZoiIiHd3d2ZmZnd3d2ZmZmZmZmZmZlVVVWZmZlVVVWZmZlVVVWZmZnd3d3d3d2ZmZnd3d3d3d2ZmZnd3d2ZmZmZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d2ZmZnd3d2ZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVVVVVWZmZlVVVWZmZnd3d4iIiIiIiJmZmZmZmaqqqpmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiIiIiHd3d3d3d2ZmZmZmZmZmZlVVVWZmZlVVVVVVVVVVVWZmZnd3d2ZmZnd3d3d3d3d3d2ZmZnd3d2ZmZmZmZmZmZnd3d2ZmZnd3d3d3d2ZmZmZmZnd3d2ZmZnd3d3d3d2ZmZnd3d2ZmZnd3d2ZmZmZmZnd3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZlVVVWZmZmZmZmZmZoiIiJmZmaqqqqqqqpmZmaqqqqqqqqqqqqqqqoiIiGZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZlVVVURERDMzM1VVVWZmZmZmZkRERERERERERFVVVURERERERERERERERERERCIiIjMzMyIiIjMzM0RERERERDMzMzMzMyIiIjMzM4iIiMzMzLu7u6qqqqqqqqqqqpmZmZmZmYiIiIiIiIiIiGZmZlVVVURERFVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVWZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d2ZmZlVVVWZmZlVVVVVVVVVVVURERERERERERERERDMzM1VVVWZmZkRERERERERERFVVVVVVVVVVVURERERERERERERERERERFVVVVVVVURERDMzM0RERERERERERERERERERFVVVVVVVWZmZlVVVURERDMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVVVVVURERFVVVVVVVWZmZnd3d3d3d2ZmZmZmZnd3d3d3d2ZmZlVVVWZmZlVVVVVVVVVVVURERFVVVVVVVURERERERERERERERFVVVVVVVWZmZnd3d4iIiIiIiHd3d3d3d3d3d3d3d2ZmZnd3d3d3d4iIiHd3d3d3d2ZmZnd3d3d3d3d3d5mZmZmZmZmZmYiIiIiIiHd3d4iIiIiIiHd3d3d3d3d3d2ZmZnd3d2ZmZlVVVWZmZlVVVWZmZoiIiIiIiHd3d3d3d3d3d3d3d4iIiIiIiJmZmZmZmYiIiJmZmYiIiIiIiIiIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiJmZmYiIiIiIiJmZmZmZmaqqqru7u8zMzN3d3d3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////u7u7d3d3MzMzMzMzMzMzMzMzd3d3u7u7u7u7u7u7u7u7////u7u7////u7u7MzMy7u7uZmZmZmZmIiIiIiIh3d3eIiIiZmZmZmZm7u7u7u7u7u7u7u7u7u7uqqqq7u7u7u7vMzMzMzMy7u7vMzMzMzMy7u7u7u7u7u7u7u7u7u7vMzMzMzMy7u7u7u7u7u7u7u7u7u7uqqqqqqqqqqqqqqqqqqqqqqqqZmZmqqqqZmZmZmZmZmZmZmZmIiIh3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZmZmZmZmZVVVVVVVVERERERERERERERERVVVVERERERERVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3dmZmZmZmZVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIh3d3d3d3d3d3dmZmZmZmZVVVVVVVVERERERERERERVVVVERERERERVVVVmZmZERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVV3d3d3d3d3d3d3d3eIiIiIiIh3d3d3d3dmZmZVVVVmZmZVVVVmZmZmZmZ3d3dmZmZ3d3d3d3eIiIiIiIiZmZmZmZmZmZl3d3d3d3d3d3eIiIhmZmZ3d3d3d3dmZmZVVVVERERERERERERERERERERVVVVERERVVVVVVVVmZmZVVVVERERVVVVERERVVVVVVVVERERVVVV3d3eZmZnMzMzu7u7u7u7////////////u7u7////////u7u7u7u7u7u7u7u7u7u7////u7u7////u7u7////////u7u7u7u7d3d3d3d2qqqqqqqqZmZmIiIiIiIh3d3d3d3d3d3d3d3eIiIh3d3dmZmZ3d3d3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVEREQzMzMzMzMzMzNERERERERERERVVVVVVVVEREQzMzMzMzMzMzMzMzNERERERERERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZ3d3d3d3d3d3eIiIiIiIiIiIiZmZl3d3d3d3d3d3eZmZmqqqqZmZmIiIh3d3dmZmZ3d3dmZmaIiIh3d3dVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3dmZmZmZmZVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVEREQzMzNERERERERVVVVVVVVVVVVVVVVVVVVmZmZ3d3dmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVERERERERVVVVmZmaIiIiIiIiIiIiIiIiIiIiIiIiZmZmZmZm7u7uqqqqIiIhmZmZVVVVVVVVERERERERERERERERERERVVVVmZmZmZmZ3d3d3d3d3d3dmZmZ3d3d3d3dmZmZmZmZmZmaIiIiIiIhmZmZmZmZVVVVVVVVERERVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3eIiIh3d3dmZmZVVVVVVVVVVVVEREQzMzMzMzNERERERERERERVVVVVVVVmZmZmZmZmZmZ3d3dmZmZmZmZ3d3eIiIh3d3dVVVVVVVVVVVVVVVVmZmZmZmZ3d3dmZmZ3d3dmZmZVVVVVVVV3d3dmZmZ3d3d3d3eIiIiIiIh3d3dVVVVVVVVERERVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVEREREREREREQzMzMzMzMiIiIzMzNERERERERVVVVEREREREREREREREQzMzNEREREREREREQzMzNEREREREQzMzNEREQzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzNEREREREREREREREREREQzMzNEREREREQzMzMzMzMzMzNEREQzMzNEREQzMzMzMzNEREQzMzMzMzNEREQzMzMzMzMzMzNERERVVVVEREQzMzNEREQzMzNERERERERERERERERVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmaIiIiIiIh3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZ3d3d3d3d3d3dmZmZ3d3d3d3d3d3d3d3dmZmZ3d3dmZmZmZmZ3d3d3d3d3d3d3d3eIiIiIiIh3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIh3d3d3d3d3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3eIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3dmZmZ3d3eIiIiZmZmqqqqqqqqZmZmZmZmqqqqqqqqZmZl3d3dmZmZERERVVVVmZmZVVVVVVVVVVVVmZmZVVVUzMzNERERERER3d3dmZmYzMzMzMzNERERVVVVERERERERVVVVVVVVEREQiIiIiIiIzMzMzMzNEREREREQzMzMzMzMzMzMzMzN3d3e7u7u7u7u7u7uqqqqZmZmZmZmZmZmZmZmZmZmIiIhmZmZERERVVVVERERVVVVERERERERVVVVmZmZVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZ3d3dmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERERERVVVVVVVVVVVVEREQzMzNVVVVVVVVmZmZVVVVVVVVERERERERERERERERERERERERERERVVVVERERERERERERVVVVVVVVmZmZmZmZVVVUzMzNEREREREREREQzMzNEREQzMzMzMzMzMzNEREQzMzNERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZmZmaIiIh3d3d3d3dmZmZ3d3eIiIiIiIh3d3dmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3eIiIh3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiZmZmIiIh3d3d3d3eIiIiZmZmZmZmZmZmIiIiIiIh3d3dmZmZmZmZ3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIh3d3eIiIh3d3eIiIiIiIiZmZmqqqqZmZmIiIiIiIh3d3eIiIiZmZmZmZmqqqqZmZmqqqq7u7vMzMzd3d3u7u7u7u7u7u7////////////////////////////////////////////////////////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u////7u7u////7u7u////////7u7u7u7u7u7u3d3d3d3dzMzMzMzM3d3dzMzMu7u7zMzMzMzMzMzM3d3dzMzM3d3dzMzMzMzMu7u7u7u7qqqqqqqqqqqqu7u7u7u7u7u7zMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7qqqqqqqqqqqqqqqqu7u7u7u7u7u7u7u7u7u7qqqqqqqqmZmZiIiIiIiId3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmVVVVVVVVREREREREREREREREREREVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3d3d3d3d3ZmZmVVVVZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmiIiIiIiIiIiId3d3iIiId3d3d3d3ZmZmZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVZmZmZmZmZmZmd3d3d3d3d3d3iIiId3d3ZmZmZmZmZmZmZmZmZmZmREREVVVVZmZmVVVVZmZmd3d3d3d3d3d3ZmZmZmZmiIiIiIiIiIiImZmZmZmZmZmZiIiId3d3d3d3ZmZmZmZmZmZmVVVVVVVVREREREREREREREREVVVVVVVVVVVVREREVVVVVVVVREREREREREREVVVVVVVVZmZmd3d3d3d3qqqqzMzM7u7u////////////////////7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u////7u7u7u7u7u7u7u7u3d3du7u7mZmZd3d3d3d3ZmZmd3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmVVVVZmZmd3d3ZmZmd3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiImZmZiIiIZmZmd3d3ZmZmVVVVVVVVVVVVVVVVREREVVVVREREVVVVREREZmZmVVVVREREREREREREREREREREREREVVVVVVVVREREREREREREREREVVVVVVVVZmZmZmZmVVVVVVVVREREVVVVVVVVVVVVZmZmZmZmd3d3ZmZmd3d3d3d3ZmZmd3d3d3d3iIiId3d3d3d3d3d3iIiId3d3ZmZmZmZmZmZmVVVVZmZmd3d3ZmZmZmZmVVVVREREREREVVVVVVVVZmZmZmZmZmZmd3d3ZmZmVVVVZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVREREREREREREVVVVVVVVVVVVVVVVZmZmZmZmVVVVREREREREREREVVVVZmZmZmZmVVVVVVVVVVVVREREVVVVREREZmZmd3d3iIiImZmZiIiId3d3iIiImZmZqqqqqqqqmZmZd3d3ZmZmZmZmZmZmZmZmVVVVREREVVVVREREREREREREVVVVVVVVd3d3d3d3d3d3d3d3iIiIZmZmZmZmZmZmiIiIiIiIZmZmZmZmVVVVVVVVVVVVZmZmVVVVREREVVVVZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3VVVVREREREREVVVVVVVVVVVVREREREREMzMzREREREREVVVVREREVVVVZmZmZmZmZmZmZmZmiIiIiIiId3d3VVVVREREREREREREZmZmZmZmZmZmZmZmd3d3ZmZmZmZmVVVVZmZmZmZmZmZmZmZmd3d3d3d3VVVVVVVVREREREREVVVVREREVVVVVVVVVVVVREREREREREREREREREREVVVVVVVVREREREREMzMzREREMzMzMzMzMzMzVVVVZmZmVVVVVVVVREREMzMzREREMzMzREREREREREREMzMzREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzVVVVVVVVREREREREMzMzREREREREREREREREMzMzREREMzMzMzMzREREMzMzREREREREMzMzMzMzMzMzMzMzMzMzVVVVVVVVREREVVVVREREMzMzREREMzMzREREMzMzREREREREREREREREREREVVVVREREREREVVVVREREVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVREREVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmVVVVZmZmZmZmVVVVVVVVREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmVVVVZmZmZmZmVVVVVVVVZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmd3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3iIiIiIiId3d3iIiId3d3iIiIiIiId3d3iIiIiIiId3d3iIiIiIiId3d3iIiId3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3ZmZmd3d3iIiIiIiIiIiId3d3iIiId3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmd3d3d3d3ZmZmZmZmd3d3d3d3d3d3d3d3mZmZqqqqmZmZiIiImZmZmZmZmZmZiIiId3d3ZmZmZmZmVVVVVVVVREREREREREREVVVVZmZmVVVVREREMzMzREREVVVVVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVMzMzMzMzIiIiIiIiMzMzREREREREMzMzMzMzMzMzMzMzVVVVqqqqu7u7u7u7mZmZmZmZiIiIiIiIiIiImZmZiIiIVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmd3d3ZmZmVVVVVVVVVVVVREREVVVVREREMzMzMzMzREREREREREREREREREREREREREREREREREREVVVVZmZmVVVVVVVVVVVVVVVVREREREREMzMzREREREREREREVVVVREREREREREREZmZmZmZmVVVVREREREREREREMzMzREREMzMzREREREREREREMzMzREREREREMzMzREREMzMzREREREREREREREREVVVVVVVVREREVVVVZmZmd3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiId3d3ZmZmd3d3ZmZmd3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3ZmZmZmZmVVVVVVVVZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmZmZmd3d3iIiImZmZmZmZmZmZiIiIiIiIiIiIiIiImZmZqqqqqqqqu7u7zMzM3d3d3d3d7u7u7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7v///+7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3czMzLu7u7u7u6qqqqqqqru7u6qqqszMzMzMzMzMzMzMzMzMzN3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u8zMzMzMzLu7u7u7u7u7u7u7u6qqqru7u6qqqqqqqpmZmZmZmYiIiIiIiIiIiHd3d2ZmZmZmZmZmZlVVVVVVVURERERERERERERERERERERERFVVVVVVVURERERERERERERERFVVVVVVVWZmZmZmZmZmZmZmZnd3d3d3d2ZmZnd3d2ZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d2ZmZmZmZlVVVVVVVURERFVVVWZmZnd3d2ZmZlVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVWZmZnd3d4iIiJmZmZmZmXd3d3d3d2ZmZlVVVWZmZlVVVVVVVVVVVVVVVWZmZmZmZlVVVWZmZnd3d4iIiIiIiHd3d3d3d4iIiIiIiJmZmYiIiIiIiJmZmYiIiHd3d2ZmZlVVVVVVVVVVVURERERERDMzMzMzM0RERFVVVVVVVVVVVVVVVVVVVURERERERDMzM0RERGZmZnd3d4iIiKqqqszMzN3d3e7u7v///////+7u7v///+7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7szMzIiIiGZmZlVVVVVVVURERERERDMzM0RERERERDMzM0RERERERFVVVURERERERFVVVVVVVURERERERFVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZlVVVWZmZmZmZlVVVVVVVVVVVURERFVVVVVVVVVVVURERERERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVURERFVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZmZmZlVVVVVVVWZmZnd3d3d3d2ZmZmZmZmZmZmZmZnd3d2ZmZlVVVWZmZlVVVXd3d4iIiHd3d1VVVURERERERFVVVURERGZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZnd3d4iIiHd3d2ZmZmZmZlVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVURERFVVVVVVVVVVVURERFVVVURERERERFVVVVVVVVVVVWZmZlVVVURERERERERERERERERERFVVVWZmZlVVVVVVVURERFVVVURERERERGZmZnd3d5mZmZmZmYiIiHd3d3d3d5mZmaqqqqqqqoiIiFVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVURERERERERERFVVVWZmZmZmZnd3d3d3d4iIiHd3d3d3d4iIiIiIiGZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVWZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d2ZmZmZmZkRERERERERERERERERERFVVVURERERERFVVVURERFVVVURERERERFVVVVVVVWZmZmZmZmZmZoiIiHd3d2ZmZlVVVURERERERFVVVVVVVWZmZmZmZnd3d3d3d3d3d2ZmZlVVVWZmZmZmZmZmZmZmZnd3d2ZmZkRERERERERERERERFVVVURERFVVVVVVVVVVVURERERERFVVVURERFVVVVVVVVVVVURERERERERERERERDMzM1VVVVVVVWZmZmZmZlVVVVVVVURERERERERERERERERERERERERERERERDMzM0RERERERDMzMzMzMzMzMzMzMzMzMyIiIkRERGZmZmZmZlVVVURERERERERERERERERERDMzMzMzM0RERDMzM0RERDMzM0RERDMzM0RERDMzMzMzMzMzM0RERFVVVVVVVWZmZmZmZkRERFVVVURERERERDMzM0RERERERERERERERERERERERERERERERERERERERERERERERFVVVVVVVVVVVVVVVWZmZkRERFVVVURERERERERERERERFVVVWZmZlVVVVVVVVVVVVVVVWZmZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZlVVVVVVVVVVVVVVVURERERERERERFVVVURERERERERERERERERERFVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZlVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZnd3d2ZmZnd3d3d3d3d3d2ZmZnd3d3d3d2ZmZnd3d2ZmZmZmZmZmZmZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVXd3d2ZmZlVVVVVVVWZmZmZmZlVVVWZmZnd3d3d3d3d3d3d3d3d3d3d3d4iIiKqqqqqqqqqqqoiIiJmZmZmZmYiIiIiIiHd3d2ZmZlVVVWZmZlVVVVVVVURERDMzM0RERGZmZlVVVURERDMzM1VVVWZmZkRERDMzM0RERERERERERFVVVWZmZmZmZkRERERERDMzMzMzMyIiIjMzM0RERERERERERDMzMzMzMzMzM0RERJmZmbu7u6qqqqqqqpmZmYiIiIiIiJmZmYiIiHd3d2ZmZlVVVURERFVVVVVVVVVVVURERERERERERFVVVWZmZlVVVWZmZmZmZnd3d2ZmZmZmZmZmZnd3d3d3d2ZmZlVVVURERERERFVVVURERERERERERERERERERERERERERERERERERERERERERERERFVVVWZmZlVVVURERFVVVWZmZmZmZlVVVVVVVVVVVURERFVVVURERERERERERERERERERFVVVWZmZlVVVURERERERERERDMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERDMzM0RERFVVVURERFVVVURERERERFVVVVVVVWZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZnd3d2ZmZmZmZnd3d2ZmZmZmZmZmZnd3d3d3d2ZmZnd3d2ZmZnd3d2ZmZmZmZnd3d2ZmZnd3d3d3d3d3d3d3d3d3d4iIiIiIiHd3d2ZmZnd3d2ZmZlVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZnd3d3d3d3d3d4iIiIiIiIiIiIiIiHd3d3d3d2ZmZmZmZnd3d2ZmZmZmZoiIiJmZmbu7u5mZmZmZmYiIiJmZmaqqqru7u8zMzMzMzN3d3e7u7u7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////u7u7////////u7u7u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7////u7u7////u7u7////u7u7d3d3d3d3MzMzMzMy7u7vMzMy7u7u7u7u7u7vMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMy7u7vMzMy7u7vMzMzMzMzMzMzMzMzMzMzd3d3MzMzMzMzMzMy7u7u7u7u7u7uqqqqqqqqqqqqqqqqqqqqqqqqZmZmZmZmIiIh3d3d3d3dmZmZVVVVERERERERERERERERERERVVVVERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZ3d3d3d3d3d3eIiIiIiIiIiIh3d3d3d3dmZmZVVVVmZmZVVVVVVVVVVVVERERVVVVmZmZ3d3dmZmZVVVVERERVVVVERERVVVVERERVVVVVVVVmZmZVVVVVVVVVVVVmZmZ3d3eIiIiIiIiIiIiZmZmIiIhmZmZVVVVVVVVmZmZmZmZ3d3dmZmZmZmZmZmZVVVVmZmZVVVV3d3eIiIh3d3eIiIiZmZmZmZmIiIiIiIiqqqqZmZmZmZl3d3eIiIh3d3dmZmZEREREREREREQzMzNERERERERVVVVERERVVVVmZmZVVVVVVVVVVVVERERVVVVmZmaIiIiqqqrMzMzu7u7u7u7u7u7////////u7u7////////////u7u7u7u7u7u7d3d3d3d3d3d3MzMzMzMzMzMzMzMzd3d3d3d3u7u7u7u7u7u7u7u7////u7u7d3d3d3d2qqqqZmZl3d3d3d3dVVVVERERVVVVERERERERERERVVVVVVVV3d3d3d3dmZmZVVVV3d3dmZmZmZmZmZmZmZmZmZmZ3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVERERERERERERERERERERERERERERERERVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZmZmZVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3dVVVVVVVVVVVVERERVVVVVVVVVVVVmZmZVVVVmZmZmZmZVVVVmZmZmZmZmZmaIiIh3d3dmZmZmZmZVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZVVVVmZmZERERERERVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVERERERERVVVVVVVVERERVVVVmZmZVVVVEREREREQzMzNERERERERERERVVVVVVVVVVVVVVVVERERERERERERERERVVVVmZmZ3d3d3d3eIiIiIiIiqqqqZmZmIiIiIiIh3d3dVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVmZmZmZmZ3d3d3d3eIiIiIiIh3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZVVVVmZmZmZmZmZmZVVVVmZmZmZmZ3d3d3d3d3d3d3d3dmZmZVVVVERERERERERERERERERERVVVVVVVVVVVVmZmZVVVVERERERERERERVVVVmZmZ3d3d3d3eIiIhmZmZVVVVERERERERVVVVVVVVVVVVVVVVmZmZ3d3d3d3d3d3dmZmZVVVVVVVVmZmZ3d3dmZmZVVVVVVVVERERERERERERERERERERVVVVERERVVVVERERVVVVVVVVVVVVERERERERERERVVVVERERVVVVEREQzMzNERERERERVVVVVVVVERERVVVVVVVVVVVVVVVVERERVVVUzMzMzMzNEREQzMzMzMzNEREQzMzNEREQzMzMzMzMzMzMzMzNERERERERmZmZVVVVEREREREREREREREREREQzMzNEREQzMzNEREREREQzMzNEREQzMzNEREQzMzNERERERERERERVVVVmZmZVVVVVVVVEREREREREREREREREREREREQzMzMzMzNERERERERERERERERERERERERERERERERERERVVVVVVVVVVVVVVVVEREREREREREREREQzMzNEREQzMzMzMzNERERmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVERERVVVVVVVVVVVVERERVVVVERERVVVVVVVVERERVVVVVVVVERERERERVVVVERERVVVVVVVVmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZmZmZ3d3dmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVV3d3dmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3dVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVmZmZmZmZmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZ3d3d3d3dmZmZ3d3d3d3d3d3eIiIiIiIh3d3eIiIh3d3d3d3d3d3dmZmZmZmZmZmZVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZ3d3dmZmZ3d3dmZmZ3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3eIiIh3d3eIiIh3d3dmZmZ3d3eIiIiZmZm7u7u7u7uqqqqZmZmIiIiZmZmIiIh3d3eIiIhmZmZVVVVmZmZVVVVVVVVEREQzMzMzMzNERERVVVVERERERERVVVVmZmZVVVVEREQzMzNERERERERmZmZ3d3dmZmZVVVVEREREREQzMzMiIiIzMzNEREREREQzMzMzMzMzMzNEREQzMzNmZmaqqqqqqqqqqqqZmZmIiIh3d3d3d3eIiIh3d3dmZmZVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dVVVVVVVVEREREREREREREREREREQzMzNEREREREREREREREREREQzMzNERERERERERERVVVVVVVVERERERERmZmZ3d3dmZmZmZmZmZmZVVVVVVVVERERERERERERVVVVERERERERVVVVmZmZEREREREREREREREQzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREREREREREREREQzMzNEREQzMzNERERERERVVVVVVVVmZmZmZmZmZmZERERVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZ3d3eIiIiIiIiZmZmIiIiIiIh3d3d3d3d3d3dmZmZ3d3d3d3d3d3d3d3eIiIiZmZmqqqqqqqqZmZmqqqqqqqq7u7vd3d3d3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u7u7u////////7u7u////////////////////7u7u////7u7u3d3d3d3d3d3dzMzMzMzMu7u7zMzMzMzMzMzMzMzM3d3dzMzM3d3du7u7u7u7qqqqu7u7u7u7u7u7zMzMzMzMzMzMzMzMzMzM3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMu7u7u7u7qqqqu7u7qqqqmZmZqqqqqqqqmZmZmZmZd3d3d3d3VVVVVVVVREREREREMzMzREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmd3d3d3d3iIiIiIiIiIiId3d3d3d3d3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmd3d3iIiId3d3iIiId3d3d3d3ZmZmd3d3ZmZmVVVVZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmVVVVZmZmiIiImZmZiIiImZmZqqqqu7u7mZmZmZmZmZmZmZmZiIiIZmZmVVVVVVVVVVVVREREVVVVREREREREVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVZmZmiIiIqqqqzMzM3d3d////////////////////7u7u////7u7u////7u7u7u7u7u7u3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzM3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3dzMzMu7u7mZmZiIiIiIiId3d3d3d3ZmZmVVVVZmZmd3d3ZmZmiIiImZmZd3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3VVVVREREVVVVREREVVVVVVVVREREREREREREREREREREREREMzMzREREREREREREMzMzREREMzMzREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3iIiId3d3iIiIiIiId3d3d3d3ZmZmZmZmZmZmZmZmZmZmd3d3ZmZmVVVVVVVVVVVVZmZmZmZmd3d3d3d3ZmZmd3d3ZmZmZmZmd3d3VVVVZmZmZmZmZmZmZmZmd3d3ZmZmZmZmVVVVZmZmZmZmZmZmVVVVVVVVZmZmZmZmd3d3ZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmiIiIiIiIZmZmVVVVVVVVVVVVVVVVREREREREREREREREVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREVVVVREREVVVVVVVVVVVVZmZmVVVVREREMzMzREREREREREREREREVVVVVVVVVVVVVVVVVVVVREREREREREREREREVVVVREREZmZmiIiImZmZqqqqiIiId3d3d3d3VVVVREREREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmZmZmd3d3d3d3d3d3iIiId3d3VVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVZmZmd3d3d3d3d3d3d3d3ZmZmVVVVREREREREREREREREREREVVVVVVVVVVVVVVVVZmZmZmZmVVVVREREVVVVVVVVd3d3d3d3ZmZmZmZmZmZmVVVVMzMzREREREREVVVVVVVVVVVVVVVVZmZmd3d3ZmZmVVVVVVVVVVVVZmZmZmZmVVVVREREVVVVREREREREMzMzREREREREREREREREREREREREVVVVVVVVVVVVVVVVREREREREREREVVVVREREREREREREREREREREREREMzMzREREREREVVVVVVVVVVVVVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREMzMzMzMzREREREREREREMzMzREREMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzREREREREVVVVZmZmVVVVREREREREREREMzMzMzMzREREMzMzREREREREMzMzMzMzREREMzMzREREREREREREREREREREVVVVVVVVVVVVVVVVREREVVVVREREREREREREREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVREREVVVVVVVVREREVVVVREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmiIiId3d3ZmZmVVVVZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVZmZmVVVVVVVVZmZmd3d3d3d3ZmZmd3d3d3d3ZmZmVVVVVVVVZmZmZmZmd3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3ZmZmd3d3d3d3d3d3d3d3iIiIiIiImZmZmZmZqqqqmZmZmZmZiIiIiIiIiIiImZmZiIiId3d3d3d3d3d3d3d3d3d3ZmZmZmZmd3d3ZmZmd3d3ZmZmd3d3d3d3ZmZmd3d3ZmZmd3d3ZmZmZmZmd3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3d3d3mZmZu7u7qqqqqqqqqqqqmZmZiIiIiIiIiIiIiIiId3d3ZmZmVVVVVVVVVVVVREREREREREREVVVVREREREREREREREREZmZmZmZmREREMzMzREREVVVVVVVVVVVVd3d3d3d3VVVVMzMzMzMzMzMzIiIiIiIiMzMzREREREREMzMzMzMzMzMzREREREREiIiIu7u7qqqqmZmZmZmZiIiId3d3d3d3d3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVd3d3ZmZmZmZmVVVVVVVVZmZmZmZmZmZmd3d3ZmZmZmZmVVVVREREREREREREREREMzMzREREREREREREREREREREMzMzMzMzMzMzREREREREREREVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVREREREREVVVVVVVVVVVVREREVVVVVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREREREMzMzREREMzMzMzMzREREREREREREREREVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVREREVVVVREREVVVVVVVVVVVVREREREREREREVVVVREREREREVVVVREREVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3iIiIiIiIiIiIiIiId3d3d3d3ZmZmd3d3d3d3d3d3d3d3iIiImZmZmZmZqqqqqqqqu7u7u7u7u7u73d3d3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3czMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u6qqqqqqqru7u7u7u8zMzMzMzMzMzN3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u6qqqru7u6qqqqqqqqqqqoiIiIiIiHd3d2ZmZlVVVVVVVURERFVVVURERERERFVVVVVVVVVVVVVVVVVVVWZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d4iIiIiIiHd3d3d3d2ZmZlVVVVVVVVVVVURERFVVVURERFVVVURERFVVVVVVVURERERERFVVVVVVVVVVVWZmZmZmZlVVVVVVVWZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZlVVVVVVVVVVVVVVVWZmZlVVVWZmZnd3d3d3d2ZmZmZmZnd3d3d3d2ZmZmZmZnd3d5mZmbu7u6qqqpmZmZmZmZmZmZmZmYiIiHd3d3d3d2ZmZlVVVVVVVURERFVVVVVVVWZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZoiIiJmZmczMzO7u7u7u7v///////+7u7u7u7v///////+7u7u7u7v///+7u7u7u7u7u7u7u7szMzN3d3d3d3d3d3d3d3d3d3d3d3e7u7t3d3e7u7t3d3d3d3e7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7szMzKqqqoiIiHd3d3d3d3d3d3d3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVURERERERERERDMzM0RERDMzMzMzMzMzM0RERDMzMzMzMzMzM0RERDMzM1VVVURERERERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d2ZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZkRERFVVVXd3d4iIiGZmZmZmZoiIiHd3d2ZmZmZmZnd3d3d3d3d3d3d3d2ZmZnd3d2ZmZmZmZmZmZnd3d2ZmZmZmZmZmZnd3d3d3d1VVVVVVVURERFVVVXd3d3d3d3d3d3d3d3d3d3d3d2ZmZlVVVWZmZlVVVVVVVVVVVVVVVURERFVVVURERFVVVVVVVURERERERFVVVVVVVVVVVVVVVWZmZkRERERERERERFVVVVVVVVVVVURERFVVVURERERERFVVVURERERERFVVVURERERERERERERERFVVVVVVVVVVVURERDMzM0RERERERERERERERERERERERERERFVVVVVVVURERERERERERERERERERERERFVVVXd3d4iIiHd3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZnd3d3d3d3d3d2ZmZmZmZlVVVVVVVURERFVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d4iIiHd3d3d3d1VVVVVVVVVVVURERERERERERERERERERFVVVURERFVVVVVVVVVVVVVVVURERFVVVURERFVVVXd3d2ZmZmZmZmZmZlVVVURERERERERERERERFVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVWZmZmZmZkRERERERERERERERERERDMzMzMzM0RERERERERERERERERERFVVVVVVVVVVVURERERERERERFVVVURERERERERERERERFVVVURERERERERERERERERERERERFVVVURERFVVVURERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERDMzM0RERDMzMzMzM0RERERERERERERERERERERERDMzMzMzM0RERDMzM0RERDMzMzMzM0RERERERERERFVVVURERERERERERERERDMzM0RERERERDMzMzMzMzMzM0RERERERDMzMzMzM0RERDMzMzMzM0RERERERFVVVVVVVVVVVURERERERERERFVVVWZmZkRERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVVVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZmZmZnd3d2ZmZnd3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d3d3d2ZmZnd3d2ZmZmZmZmZmZnd3d2ZmZnd3d2ZmZnd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiKqqqqqqqqqqqqqqqpmZmYiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d4iIiJmZmaqqqru7u6qqqqqqqpmZmZmZmZmZmZmZmYiIiHd3d3d3d2ZmZlVVVURERERERERERFVVVVVVVVVVVURERERERERERFVVVWZmZmZmZkRERDMzM1VVVWZmZlVVVVVVVWZmZmZmZkRERERERDMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzM0RERFVVVZmZmaqqqqqqqqqqqpmZmYiIiHd3d3d3d3d3d3d3d2ZmZlVVVVVVVVVVVVVVVURERFVVVVVVVWZmZmZmZmZmZlVVVWZmZmZmZnd3d3d3d2ZmZnd3d3d3d2ZmZkRERFVVVVVVVURERERERERERDMzM0RERERERERERERERDMzM0RERERERERERFVVVWZmZlVVVVVVVVVVVWZmZlVVVVVVVVVVVURERERERERERERERFVVVURERFVVVURERERERERERFVVVVVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERDMzMzMzM0RERERERERERERERERERERERERERERERERERERERERERERERFVVVURERERERERERERERERERERERFVVVURERFVVVURERERERERERERERERERERERERERERERFVVVURERERERERERFVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERERERFVVVVVVVWZmZmZmZnd3d3d3d4iIiIiIiIiIiHd3d2ZmZmZmZmZmZoiIiHd3d2ZmZnd3d4iIiJmZmaqqqru7u7u7u7u7u8zMzMzMzO7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7u7u7d3d3u7u7u7u7d3d3d3d3u7u7d3d3d3d3d3d3MzMzMzMzMzMy7u7uqqqqqqqqZmZmqqqqqqqq7u7u7u7u7u7vMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7vMzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7uqqqq7u7uqqqqqqqqqqqqZmZmIiIh3d3dmZmZmZmZmZmZVVVVmZmZVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVmZmZ3d3dmZmZ3d3d3d3d3d3d3d3dmZmZ3d3eIiIiIiIh3d3d3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVERERVVVVERERERERVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZ3d3d3d3d3d3dmZmZmZmZmZmZVVVVERERVVVVVVVVVVVVVVVVmZmZVVVVVVVVmZmZ3d3d3d3dmZmaIiIiIiIiIiIh3d3d3d3eZmZmZmZmqqqqqqqqZmZmIiIh3d3d3d3dmZmZVVVVVVVVERERERERERERERERVVVVmZmZmZmZ3d3d3d3d3d3d3d3dmZmZmZmZmZmaZmZnMzMzu7u7u7u7////////////////////////////////////u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3u7u7d3d3d3d3d3d3d3d3u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3MzMyqqqpmZmZVVVVVVVVVVVVVVVVVVVVVVVVEREREREREREREREREREQzMzNERERERERERERERERERERERERERERVVVVmZmZmZmZ3d3dVVVVVVVVEREQzMzMzMzMzMzNERERVVVVEREQzMzMzMzNEREREREQzMzNVVVVEREREREREREQzMzMzMzNEREREREQzMzMzMzNEREREREQzMzNERERERERERERVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVVERERVVVVmZmZ3d3dVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZVVVVmZmZ3d3d3d3dmZmZmZmZmZmZVVVVVVVVVVVVmZmZmZmZ3d3d3d3dmZmZ3d3dmZmZmZmZmZmZVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVmZmZVVVVERERERERVVVVVVVVERERERERERERERERERERVVVVVVVVVVVVERERVVVVVVVVERERERERVVVVERERmZmZVVVVEREREREREREREREQzMzNERERERERERERERERVVVVERERERERERERERERVVVVVVVVERERVVVVmZmZ3d3d3d3dmZmZVVVVERERVVVVERERERERERERERERVVVVmZmZmZmZVVVVVVVVERERVVVVVVVVmZmZmZmZ3d3eIiIh3d3d3d3dmZmZmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVVVVVmZmZmZmaIiIh3d3d3d3dmZmZmZmZEREREREREREREREREREREREQzMzNERERVVVVVVVVVVVVERERVVVVERERVVVVVVVVmZmZ3d3dmZmZmZmZVVVVEREQzMzNERERERERVVVVVVVVVVVVVVVVERERVVVVERERERERERERVVVVmZmZmZmZVVVVEREREREREREREREREREREREREREQzMzNERERVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERERERVVVVEREREREQzMzMzMzNERERVVVVVVVVEREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREQzMzMzMzMzMzNEREQzMzNEREREREREREREREREREQzMzMzMzMzMzMzMzNEREREREQzMzNEREREREREREREREREREREREREREREREQzMzNEREQzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzNERERERERERERmZmZmZmZVVVVERERVVVVVVVVVVVVERERERERERERVVVVmZmZVVVVmZmZ3d3dERERVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZVVVVmZmZmZmZVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3dmZmZmZmZ3d3d3d3d3d3dmZmZ3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3dmZmZmZmZ3d3dmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3eIiIiIiIiIiIiIiIiZmZmIiIiIiIiIiIiZmZmZmZmZmZmqqqqZmZmZmZmIiIiIiIiIiIiIiIh3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3eIiIiqqqqqqqq7u7uqqqqZmZmZmZmZmZmZmZmIiIiIiIh3d3dmZmZVVVVVVVVERERERERERERERERmZmZVVVUzMzNVVVVERERVVVVVVVVmZmZERERERERmZmZVVVVERERERERVVVVmZmZEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzNERERERERERER3d3eZmZmqqqqqqqqqqqqZmZmIiIiIiIiIiIh3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZ3d3d3d3d3d3dmZmZmZmZmZmZVVVVVVVVVVVVEREREREREREREREREREREREREREREREREREREREQzMzNERERERERERERVVVVmZmZmZmZVVVVVVVVVVVVERERERERERERERERERERVVVVVVVVVVVVERERERERVVVVVVVVVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzNEREREREREREQzMzNERERERERVVVVERERERERVVVVERERERERERERERERERERERERERERVVVVERERERERERERERERVVVVVVVVERERERERERERERERERERERERERERERERERERERERERERVVVVVVVVmZmZERERERERERERERERVVVVVVVVERERVVVVERERVVVVVVVVERERVVVVVVVVmZmZ3d3eIiIiIiIiZmZmZmZl3d3dmZmZmZmZ3d3eIiIiZmZmIiIh3d3d3d3eIiIiqqqq7u7u7u7u7u7vMzMzMzMzu7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMu7u7qqqqqqqqqqqqu7u7u7u7zMzMu7u7zMzMzMzMzMzMu7u7zMzMu7u7zMzMzMzMzMzMzMzMzMzMzMzM3d3dzMzMzMzMzMzMzMzMu7u7zMzMu7u7qqqqu7u7qqqqqqqqu7u7qqqqqqqqmZmZiIiIiIiId3d3ZmZmZmZmd3d3d3d3ZmZmZmZmZmZmd3d3d3d3d3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiIiIiId3d3d3d3d3d3ZmZmZmZmVVVVZmZmZmZmVVVVZmZmZmZmVVVVREREREREREREREREREREVVVVVVVVVVVVZmZmVVVVd3d3d3d3ZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmVVVVVVVVVVVVREREREREVVVVVVVVVVVVZmZmd3d3ZmZmd3d3d3d3iIiIiIiId3d3d3d3d3d3iIiIiIiImZmZmZmZmZmZd3d3d3d3ZmZmZmZmZmZmVVVVVVVVREREREREVVVVVVVVZmZmd3d3iIiIiIiIiIiImZmZmZmZmZmZmZmZu7u7zMzM7u7u////////////////////7u7u////////////7u7u7u7u7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3dzMzMzMzM3d3d7u7u7u7u7u7u7u7u7u7u////7u7u7u7u7u7u3d3d7u7u3d3du7u7mZmZiIiIZmZmVVVVVVVVREREREREREREVVVVVVVVVVVVVVVVREREREREREREREREMzMzMzMzREREVVVVZmZmmZmZu7u7qqqqiIiId3d3VVVVVVVVREREMzMzREREVVVVREREMzMzIiIiMzMzMzMzMzMzMzMzREREREREREREMzMzREREMzMzREREMzMzREREREREREREREREMzMzREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVZmZmVVVVZmZmZmZmd3d3d3d3iIiId3d3d3d3d3d3ZmZmVVVVVVVVZmZmZmZmZmZmVVVVVVVVREREVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVZmZmVVVVREREREREVVVVREREVVVVVVVVREREREREREREREREVVVVVVVVVVVVVVVVREREVVVVREREREREREREVVVVREREMzMzREREMzMzREREREREREREREREREREREREREREVVVVREREVVVVVVVVVVVVVVVVREREVVVVZmZmZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVVVVVREREREREVVVVZmZmd3d3iIiIiIiId3d3d3d3VVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREVVVVZmZmd3d3d3d3d3d3ZmZmVVVVREREREREREREREREMzMzREREREREREREREREVVVVREREREREMzMzREREREREVVVVZmZmd3d3VVVVZmZmREREREREMzMzREREREREVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREZmZmZmZmVVVVREREREREREREREREMzMzREREREREREREREREVVVVZmZmVVVVVVVVREREMzMzREREVVVVVVVVVVVVREREMzMzREREREREREREREREREREMzMzREREMzMzREREVVVVREREMzMzMzMzREREREREREREREREMzMzIiIiMzMzMzMzREREMzMzMzMzMzMzREREREREREREMzMzMzMzREREREREMzMzREREREREREREMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREVVVVREREMzMzMzMzREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzREREREREVVVVVVVVREREVVVVREREVVVVREREMzMzREREREREREREd3d3ZmZmZmZmZmZmZmZmVVVVREREVVVVZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiId3d3iIiId3d3d3d3d3d3d3d3d3d3iIiIZmZmd3d3d3d3d3d3d3d3iIiId3d3iIiIiIiId3d3d3d3iIiId3d3d3d3iIiId3d3iIiId3d3iIiIiIiIiIiIiIiImZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3iIiId3d3d3d3d3d3ZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmVVVVZmZmZmZmVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3iIiIZmZmiIiImZmZqqqqqqqqmZmZmZmZmZmZqqqqmZmZiIiId3d3ZmZmZmZmVVVVVVVVVVVVREREVVVVZmZmVVVVREREREREZmZmVVVVREREVVVVVVVVVVVVVVVVZmZmVVVVMzMzMzMzVVVVZmZmVVVVREREREREMzMzMzMzIiIiMzMzMzMzREREMzMzIiIiMzMzMzMzREREREREVVVVd3d3mZmZu7u7qqqqqqqqiIiIiIiIiIiId3d3d3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmVVVVVVVVREREREREREREREREVVVVREREREREREREREREREREREREREREVVVVVVVVZmZmZmZmZmZmZmZmVVVVVVVVREREVVVVREREVVVVVVVVREREVVVVVVVVREREVVVVZmZmVVVVVVVVVVVVMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzREREMzMzREREREREREREREREREREREREVVVVREREREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVREREREREREREREREREREREREREREREREVVVVREREREREVVVVVVVVVVVVVVVVREREREREREREVVVVREREREREVVVVREREVVVVVVVVVVVVVVVVZmZmd3d3iIiIiIiIiIiIiIiId3d3d3d3ZmZmZmZmiIiImZmZqqqqmZmZiIiImZmZmZmZu7u7u7u7zMzM3d3d3d3d3d3d////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u7u7u8zMzLu7u8zMzMzMzMzMzN3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u8zMzLu7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqpmZmYiIiJmZmYiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZnd3d2ZmZnd3d2ZmZnd3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d2ZmZmZmZlVVVVVVVURERFVVVVVVVVVVVVVVVVVVVURERERERFVVVURERFVVVWZmZlVVVVVVVVVVVVVVVWZmZmZmZnd3d3d3d3d3d4iIiHd3d4iIiIiIiHd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZlVVVURERFVVVVVVVVVVVWZmZnd3d2ZmZnd3d4iIiIiIiIiIiIiIiHd3d3d3d4iIiIiIiIiIiIiIiIiIiGZmZnd3d2ZmZmZmZmZmZlVVVWZmZlVVVVVVVXd3d3d3d3d3d3d3d5mZmaqqqqqqqru7u8zMzN3d3d3d3e7u7v///////////////////////////////////////////////////////+7u7v///+7u7v///+7u7v///////+7u7v///+7u7t3d3czMzLu7u7u7u8zMzMzMzN3d3e7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3czMzLu7u5mZmXd3d2ZmZmZmZmZmZlVVVWZmZnd3d4iIiHd3d3d3d2ZmZmZmZkRERERERERERFVVVVVVVXd3d6qqqqqqqpmZmYiIiGZmZmZmZmZmZkRERERERDMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzM0RERERERERERERERERERERERDMzM0RERERERERERERERFVVVVVVVURERERERDMzM0RERDMzM0RERERERFVVVURERFVVVURERFVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZmZmZmZmZlVVVXd3d4iIiIiIiIiIiJmZmYiIiHd3d3d3d2ZmZlVVVWZmZmZmZmZmZkRERERERERERFVVVURERFVVVVVVVWZmZlVVVVVVVURERFVVVVVVVURERFVVVVVVVURERFVVVVVVVVVVVVVVVVVVVURERFVVVWZmZlVVVVVVVURERERERERERFVVVURERFVVVURERFVVVURERFVVVVVVVVVVVURERFVVVVVVVVVVVURERFVVVVVVVURERERERDMzM0RERDMzM0RERERERERERERERERERERERERERERERERERERERERERFVVVURERERERERERFVVVVVVVURERERERFVVVURERFVVVURERERERERERERERERERERERERERERERERERERERERERFVVVXd3d3d3d3d3d3d3d2ZmZkRERFVVVURERFVVVURERERERFVVVURERFVVVWZmZlVVVVVVVURERERERERERERERFVVVWZmZmZmZnd3d3d3d2ZmZkRERDMzM0RERDMzM0RERDMzM0RERDMzM0RERERERERERERERERERERERDMzM0RERERERGZmZnd3d2ZmZlVVVURERDMzMzMzM0RERERERFVVVVVVVVVVVVVVVVVVVTMzM0RERERERERERFVVVVVVVWZmZkRERERERERERERERERERERERERERERERERERERERFVVVVVVVURERERERDMzMzMzMzMzM0RERFVVVVVVVVVVVURERDMzM0RERERERERERDMzM0RERDMzM0RERERERDMzM0RERERERDMzMzMzMzMzM1VVVURERERERDMzMzMzM0RERERERERERDMzMzMzM0RERERERDMzMzMzM0RERDMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERDMzM0RERERERDMzM0RERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERFVVVVVVVURERERERFVVVVVVVURERDMzM0RERERERERERGZmZlVVVWZmZlVVVXd3d2ZmZmZmZmZmZnd3d5mZmYiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d3d3d2ZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZlVVVWZmZlVVVWZmZlVVVWZmZmZmZlVVVWZmZlVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d4iIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZmZmZnd3d2ZmZnd3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d4iIiHd3d2ZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d2ZmZnd3d3d3d4iIiHd3d3d3d3d3d3d3d3d3d4iIiHd3d2ZmZoiIiHd3d4iIiJmZmZmZmZmZmaqqqqqqqqqqqpmZmXd3d3d3d2ZmZmZmZlVVVVVVVVVVVWZmZlVVVWZmZkRERFVVVWZmZlVVVURERERERERERHd3d3d3d1VVVURERDMzMzMzM0RERFVVVURERERERERERERERERERDMzMzMzMzMzM0RERERERCIiIjMzMzMzMzMzM0RERDMzM1VVVYiIiKqqqqqqqqqqqqqqqoiIiIiIiIiIiHd3d3d3d2ZmZlVVVVVVVVVVVWZmZmZmZmZmZlVVVWZmZlVVVWZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZlVVVURERERERERERFVVVURERERERFVVVURERERERERERDMzM0RERERERFVVVVVVVVVVVWZmZlVVVVVVVVVVVURERFVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVURERFVVVVVVVVVVVURERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERDMzM0RERDMzMzMzM0RERDMzM0RERERERERERERERERERERERERERERERERERDMzM0RERERERERERERERERERERERERERFVVVVVVVURERERERERERFVVVVVVVURERFVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVXd3d4iIiIiIiIiIiHd3d3d3d2ZmZmZmZnd3d5mZmZmZmaqqqpmZmZmZmaqqqqqqqru7u7u7u8zMzMzMzN3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7////u7u7////u7u7////u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7u7u7d3d3d3d3d3d3MzMzMzMy7u7u7u7u7u7u7u7uqqqq7u7u7u7u7u7u7u7vMzMzMzMzMzMzMzMzd3d3MzMzMzMzMzMy7u7u7u7u7u7vMzMzMzMzMzMy7u7vMzMzMzMzMzMzMzMy7u7vMzMy7u7u7u7u7u7u7u7uqqqqqqqqqqqqZmZmZmZmZmZmIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3d3d3eIiIiIiIiIiIiIiIiZmZmIiIiIiIiIiIiIiIh3d3d3d3dmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZ3d3d3d3eIiIiIiIh3d3d3d3d3d3dmZmZmZmZ3d3d3d3d3d3d3d3dVVVVVVVVVVVVmZmZVVVVmZmZmZmZ3d3d3d3d3d3d3d3eIiIiZmZmIiIiIiIiIiIiIiIh3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZ3d3d3d3eIiIiIiIiZmZmqqqq7u7vMzMzd3d3u7u7u7u7////////////////////////////////////////////////////////////////////////////////////u7u7////////////////u7u7MzMy7u7u7u7vMzMzMzMzd3d3d3d3d3d3u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7d3d3u7u7d3d3d3d3MzMzMzMyqqqqZmZmZmZmZmZmqqqqqqqq7u7u7u7u7u7u7u7u7u7uqqqqZmZl3d3dmZmZmZmZVVVVmZmZmZmZmZmZ3d3dmZmZVVVVEREREREQzMzMzMzMzMzMiIiIzMzMzMzMiIiIiIiIzMzMzMzNERERVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVERERVVVVmZmZEREREREREREREREQzMzMzMzNERERERERERERERERERERVVVVVVVVmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVmZmZVVVVmZmZ3d3dmZmZmZmZmZmZ3d3eIiIiZmZmIiIh3d3eIiIiIiIhmZmZmZmZmZmZmZmZVVVVmZmZmZmZVVVVVVVVERERVVVVVVVVmZmZVVVVmZmZVVVVVVVVVVVVVVVVERERVVVVVVVVERERVVVVERERVVVVVVVVVVVVERERERERVVVVmZmZmZmZVVVVERERVVVVERERERERVVVVERERVVVVERERVVVVERERVVVVERERERERVVVVVVVVVVVVERERVVVVVVVVVVVUzMzNEREQzMzNERERERERERERVVVVEREREREREREREREREREREREREREREREREREREREQzMzNERERERERVVVVERERVVVVERERVVVVERERERERERERERERERERERERVVVVERERERERERERERERERERVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVERERERERVVVVERERERERERERERERVVVVVVVVERERERERVVVVVVVVERERERERVVVVVVVVmZmZmZmZVVVVEREQzMzMzMzNEREQzMzNEREREREQzMzNEREQzMzNEREREREREREQzMzNEREQzMzNERERmZmZ3d3dVVVVVVVVEREREREREREREREREREREREREREREREREREREREREREQzMzMzMzNERERERERmZmZVVVVVVVUzMzNEREQzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREQzMzMiIiIzMzMiIiIzMzNERERERERVVVVVVVVERERVVVVVVVUzMzNEREQzMzNEREQzMzNEREREREREREREREREREQzMzMzMzMzMzNERERERERERERERERVVVVVVVVEREQzMzMzMzNEREREREQzMzNEREQzMzNEREQzMzNEREREREQzMzMzMzMiIiIiIiIzMzMzMzMzMzNEREQzMzNVVVVVVVVEREQiIiIzMzNEREQzMzNEREREREQzMzMzMzNEREQzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzNERERVVVVVVVVERERERERVVVVVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmaIiIiIiIiIiIh3d3eIiIiZmZmIiIiIiIiIiIh3d3d3d3d3d3d3d3dmZmZmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZVVVVVVVVmZmZVVVVmZmZmZmZVVVVmZmZVVVVmZmZmZmZmZmZVVVVmZmZmZmZmZmZ3d3dmZmZVVVVmZmZmZmZmZmZVVVVmZmZmZmZmZmZVVVVmZmZ3d3dmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZ3d3eIiIiZmZmIiIiIiIiIiIiIiIh3d3eIiIiIiIh3d3dmZmZ3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3d3d3eIiIh3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3d3d3d3d3dmZmZ3d3dmZmZmZmZ3d3d3d3dmZmZ3d3d3d3eIiIiZmZmqqqqqqqqqqqqZmZmZmZmIiIiIiIh3d3d3d3d3d3dVVVVVVVVVVVVVVVVVVVVVVVVERERmZmZmZmZVVVVERERERERVVVVmZmZmZmZVVVUzMzNEREQzMzNERERVVVVEREQzMzNEREREREREREQzMzNEREREREREREQzMzMiIiIzMzMzMzMzMzMzMzNERERERERVVVWZmZmqqqqqqqqqqqqqqqqIiIiIiIh3d3d3d3d3d3dmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZ3d3d3d3d3d3dmZmZmZmZVVVVERERERERERERERERERERERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVERERVVVVVVVVVVVVVVVVVVVVEREQzMzNEREQzMzMzMzMiIiIzMzMzMzNEREREREREREQzMzNEREREREQzMzNEREREREREREREREQzMzNERERERERERERERERERERERERERERERERERERERERERERERERVVVVERERERERERERERERERERERERERERVVVVVVVVERERVVVVERERVVVVERERERERVVVVERERERERERERVVVVERERVVVVVVVVmZmZmZmZmZmaIiIiIiIiIiIh3d3dmZmZmZmZmZmZ3d3eIiIiZmZmZmZmqqqqqqqqZmZmqqqqqqqq7u7u7u7vMzMzd3d3u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u3d3d7u7u3d3d3d3d3d3d3d3dzMzMzMzMzMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7zMzMzMzM3d3d3d3d3d3dzMzMzMzMu7u7u7u7u7u7u7u7qqqqqqqqqqqqqqqqu7u7u7u7zMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqqqqqmZmZiIiId3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmd3d3iIiImZmZmZmZmZmZiIiIiIiIiIiIiIiIiIiId3d3ZmZmVVVVVVVVREREVVVVREREVVVVREREREREREREVVVVVVVVZmZmZmZmZmZmd3d3ZmZmVVVVZmZmZmZmZmZmZmZmd3d3d3d3iIiId3d3iIiId3d3d3d3ZmZmZmZmd3d3ZmZmZmZmd3d3d3d3d3d3d3d3ZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3iIiIiIiImZmZmZmZiIiId3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiImZmZmZmZqqqqu7u7zMzMzMzM7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u////////////////7u7u////zMzMqqqqqqqqzMzM3d3d3d3d3d3d3d3d3d3d7u7u3d3d7u7u7u7u3d3d3d3d7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzM3d3d3d3dzMzMzMzMu7u7zMzMu7u7u7u7qqqqd3d3d3d3ZmZmVVVVZmZmZmZmVVVVVVVVREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVREREREREREREMzMzMzMzREREMzMzMzMzREREREREREREREREREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3d3d3iIiIZmZmd3d3iIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmd3d3ZmZmVVVVVVVVVVVVZmZmVVVVVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVREREVVVVREREREREREREREREVVVVVVVVREREREREVVVVVVVVVVVVZmZmVVVVVVVVREREREREREREVVVVVVVVVVVVREREVVVVREREVVVVREREREREVVVVVVVVVVVVVVVVREREVVVVVVVVREREREREMzMzREREREREREREREREREREREREREREREREVVVVREREREREREREREREREREREREMzMzREREVVVVVVVVMzMzREREREREREREVVVVREREREREVVVVREREVVVVREREVVVVREREVVVVVVVVREREREREVVVVVVVVZmZmVVVVVVVVREREREREREREREREREREREREVVVVREREVVVVVVVVREREREREVVVVREREREREVVVVVVVVREREVVVVZmZmZmZmVVVVREREMzMzMzMzMzMzMzMzREREMzMzREREMzMzREREREREREREREREMzMzMzMzMzMzREREZmZmZmZmZmZmVVVVREREREREREREREREREREREREREREREREREREREREREREMzMzREREMzMzREREVVVVVVVVREREMzMzREREREREREREMzMzREREMzMzMzMzMzMzREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREVVVVVVVVVVVVREREMzMzREREREREREREREREREREREREREREREREREREMzMzMzMzMzMzIiIiMzMzMzMzREREREREVVVVVVVVMzMzREREREREREREMzMzREREMzMzMzMzREREMzMzREREMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzREREREREREREMzMzMzMzMzMzMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzIiIiMzMzREREVVVVVVVVMzMzMzMzVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmd3d3iIiIiIiId3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmVVVVVVVVREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVZmZmVVVVVVVVREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmZmZmZmZmVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3iIiId3d3iIiIiIiId3d3iIiIiIiId3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmd3d3ZmZmZmZmd3d3ZmZmZmZmZmZmZmZmd3d3iIiId3d3d3d3d3d3iIiIiIiIiIiId3d3d3d3d3d3ZmZmd3d3iIiImZmZqqqqqqqqmZmZiIiImZmZiIiIiIiId3d3ZmZmZmZmVVVVVVVVVVVVZmZmVVVVVVVVZmZmVVVVREREREREVVVVZmZmZmZmREREREREMzMzREREMzMzREREVVVVVVVVMzMzREREMzMzMzMzREREREREVVVVREREMzMzMzMzIiIiMzMzMzMzMzMzMzMzREREREREd3d3qqqqqqqqqqqqqqqqmZmZiIiId3d3d3d3d3d3d3d3ZmZmZmZmVVVVZmZmZmZmVVVVZmZmd3d3d3d3d3d3d3d3ZmZmZmZmd3d3ZmZmZmZmVVVVREREREREREREREREREREVVVVREREREREREREREREREREVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmVVVVREREVVVVVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREMzMzMzMzREREREREREREMzMzREREMzMzREREREREMzMzMzMzREREREREMzMzVVVVREREREREREREVVVVVVVVREREMzMzREREMzMzREREREREVVVVVVVVREREREREVVVVREREREREVVVVREREVVVVREREVVVVREREVVVVVVVVZmZmd3d3iIiImZmZiIiId3d3ZmZmVVVVZmZmZmZmiIiIqqqqqqqqqqqqqqqqqqqqqqqqqqqqu7u73d3d3d3d3d3d////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7u7u7v///+7u7u7u7u7u7t3d3d3d3czMzMzMzMzMzMzMzMzMzLu7u8zMzMzMzN3d3d3d3czMzN3d3d3d3czMzN3d3d3d3d3d3d3d3czMzMzMzKqqqru7u6qqqru7u6qqqqqqqpmZmaqqqpmZmaqqqqqqqqqqqszMzMzMzMzMzN3d3d3d3czMzN3d3czMzMzMzLu7u8zMzLu7u7u7u7u7u6qqqru7u6qqqqqqqpmZmZmZmYiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiJmZmYiIiJmZmYiIiIiIiHd3d2ZmZmZmZmZmZlVVVVVVVVVVVURERERERERERFVVVVVVVURERFVVVVVVVWZmZmZmZnd3d3d3d2ZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZlVVVWZmZmZmZnd3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d4iIiJmZmaqqqru7u8zMzN3d3d3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7v///////+7u7u7u7t3d3d3d3d3d3bu7u8zMzN3d3d3d3d3d3e7u7t3d3e7u7u7u7u7u7t3d3d3d3d3d3czMzMzMzMzMzN3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u6qqqpmZmaqqqoiIiHd3d3d3d2ZmZmZmZmZmZlVVVVVVVURERERERERERDMzM0RERFVVVURERERERERERERERFVVVVVVVWZmZmZmZmZmZmZmZnd3d4iIiHd3d3d3d2ZmZmZmZnd3d3d3d2ZmZlVVVVVVVVVVVURERERERERERERERERERERERERERERERERERDMzMzMzM0RERERERERERFVVVURERFVVVVVVVWZmZmZmZmZmZnd3d3d3d4iIiHd3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d3d3d3d3d2ZmZmZmZlVVVWZmZmZmZlVVVWZmZmZmZlVVVURERFVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVURERERERERERERERFVVVURERERERERERFVVVURERFVVVWZmZlVVVWZmZmZmZkRERFVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVURERFVVVVVVVVVVVURERERERERERERERERERERERERERERERERERERERERERERERERERERERERERDMzMzMzM0RERFVVVVVVVVVVVTMzMzMzMzMzM0RERERERERERERERERERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVWZmZlVVVVVVVVVVVURERFVVVURERERERFVVVURERFVVVVVVVURERFVVVURERERERFVVVVVVVURERERERERERGZmZlVVVVVVVURERDMzM0RERDMzMzMzMzMzMzMzM0RERDMzMzMzM0RERERERERERERERDMzMzMzM0RERGZmZmZmZlVVVVVVVURERDMzMzMzMzMzM0RERDMzM0RERDMzM0RERERERERERERERERERERERERERERERFVVVURERDMzMzMzM0RERDMzM0RERDMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVWZmZlVVVURERERERERERERERERERERERERERERERERERERERERERDMzMzMzMzMzMyIiIiIiIjMzMzMzM0RERFVVVURERDMzM0RERDMzM0RERERERDMzM0RERDMzM0RERDMzM0RERDMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzM0RERERERERERDMzMzMzMzMzM0RERDMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzM0RERFVVVURERDMzMyIiIjMzM0RERERERFVVVURERERERERERERERFVVVVVVVVVVVVVVVURERFVVVURERERERFVVVURERERERDMzMzMzMzMzM0RERERERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZlVVVWZmZlVVVWZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZnd3d3d3d3d3d3d3d2ZmZnd3d3d3d2ZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d4iIiHd3d3d3d3d3d3d3d2ZmZmZmZmZmZnd3d3d3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d2ZmZnd3d3d3d4iIiIiIiIiIiIiIiHd3d4iIiIiIiJmZmYiIiIiIiHd3d3d3d3d3d3d3d2ZmZmZmZmZmZoiIiJmZmaqqqqqqqqqqqqqqqpmZmYiIiHd3d3d3d2ZmZlVVVVVVVWZmZnd3d2ZmZlVVVWZmZlVVVURERFVVVVVVVWZmZlVVVURERERERDMzM0RERERERFVVVWZmZkRERERERERERDMzM0RERFVVVVVVVVVVVVVVVTMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzMzMzM1VVVYiIiKqqqqqqqqqqqqqqqpmZmYiIiHd3d4iIiIiIiGZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZnd3d3d3d3d3d2ZmZnd3d2ZmZmZmZmZmZkRERERERERERFVVVVVVVURERERERERERERERERERERERFVVVWZmZlVVVVVVVVVVVVVVVVVVVXd3d1VVVVVVVVVVVURERFVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVURERFVVVURERDMzMzMzMzMzMzMzM0RERDMzMzMzM0RERERERERERERERDMzMzMzMzMzMzMzM0RERERERERERERERDMzM0RERERERERERERERERERERERDMzM0RERERERERERERERFVVVURERERERERERFVVVURERERERERERERERERERERERERERERERERERERERFVVVVVVVURERFVVVVVVVVVVVWZmZnd3d4iIiIiIiIiIiHd3d2ZmZmZmZmZmZnd3d4iIiJmZmaqqqqqqqqqqqqqqqru7u7u7u8zMzN3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzd3d3d3d3MzMzd3d3d3d3d3d3d3d3u7u7d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMyqqqqqqqqZmZmqqqqqqqq7u7uqqqq7u7uqqqqqqqq7u7u7u7u7u7vMzMzMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMy7u7vMzMzMzMy7u7u7u7u7u7uqqqqZmZmqqqqIiIiIiIiIiIiZmZmZmZmIiIiIiIiIiIiIiIiZmZmZmZmZmZmZmZmIiIh3d3d3d3d3d3d3d3dVVVVVVVVmZmZmZmZVVVVERERVVVVERERERERVVVVVVVVVVVVVVVVmZmZ3d3d3d3dmZmZ3d3d3d3d3d3dmZmZmZmZ3d3d3d3d3d3eIiIh3d3d3d3dVVVVmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZ3d3dmZmZmZmZVVVVVVVVVVVVmZmZ3d3d3d3d3d3eIiIh3d3d3d3eIiIh3d3eIiIiIiIh3d3eIiIiIiIiIiIiZmZmZmZm7u7u7u7vMzMzd3d3u7u7u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7d3d2qqqq7u7vMzMzd3d3d3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3MzMzMzMzMzMy7u7u7u7vMzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7uqqqq7u7uqqqqqqqqqqqqZmZmZmZmqqqq7u7uqqqqZmZmZmZmIiIiIiIh3d3eIiIh3d3dmZmZmZmZVVVVEREREREREREQzMzNERERERERERERERERERERERERVVVVVVVVVVVVVVVVmZmZmZmZ3d3dmZmZmZmZVVVVmZmZmZmZmZmZ3d3dmZmZVVVVVVVVEREREREREREREREREREREREREREREREREREREREREREREREREREQzMzNERERVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZmZmZmZmZ3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVV3d3d3d3d3d3d3d3d3d3dmZmZVVVVVVVVERERVVVVVVVV3d3dmZmZmZmZVVVVERERERERERERERERERERVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVmZmZmZmZVVVVERERERERVVVVERERVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZERERERERERERERERERERERERERERERERERERVVVVEREREREREREREREREREQzMzMzMzNEREREREREREREREQzMzMzMzNEREREREQzMzNERERERERVVVVERERVVVVVVVVERERVVVVVVVVVVVVVVVVERERVVVVVVVV3d3dmZmZVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVERERERERVVVVERERVVVVERERERERVVVVmZmZmZmZVVVVEREQzMzNEREQzMzNEREQzMzNEREQzMzNERERERERERERERERVVVUzMzMzMzMzMzNERERmZmZmZmZmZmZEREQzMzMzMzNEREREREQzMzNEREREREQzMzNERERVVVVEREREREREREQzMzNERERVVVVVVVVEREQzMzMzMzMzMzMzMzNEREQzMzMzMzNEREQzMzNEREQzMzMzMzNEREQzMzMzMzMzMzMiIiIzMzMzMzNERERERERVVVVVVVVEREQzMzNEREQzMzNEREREREREREREREQzMzNEREQzMzNEREQzMzMiIiIiIiIzMzMiIiIzMzNEREREREREREQzMzMzMzNEREQzMzNEREREREQzMzNEREQzMzNEREQzMzMzMzMzMzMzMzMiIiIiIiIiIiIzMzNEREQzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzNERERVVVVEREQzMzMzMzMzMzMiIiIzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERVVVVVVVVERERERERERERVVVVERERERERERERVVVVERERERERVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3dmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVmZmZVVVVmZmZVVVVmZmZmZmZmZmZVVVVmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3d3d3dmZmZ3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIh3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3dmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3eIiIh3d3d3d3d3d3eIiIh3d3d3d3d3d3eIiIh3d3eIiIh3d3d3d3d3d3dmZmZ3d3dmZmZ3d3d3d3eZmZmqqqqqqqqqqqqZmZmZmZl3d3d3d3d3d3dmZmZVVVVmZmZmZmZmZmZVVVVERERERERERERVVVVVVVVmZmZmZmZEREQzMzNEREREREQzMzNERERVVVVVVVVEREREREQzMzNERERVVVVmZmZmZmZVVVVEREREREQzMzMiIiIiIiIzMzMiIiIzMzMiIiIzMzNERERmZmaZmZm7u7uqqqqqqqqZmZmIiIiIiIh3d3d3d3d3d3d3d3dmZmZVVVVVVVVmZmZmZmZVVVV3d3d3d3dmZmZVVVVmZmZ3d3dmZmZVVVVERERERERVVVVERERVVVVERERVVVVEREQzMzNERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZERERVVVVERERVVVVmZmZmZmZmZmZmZmZVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVUzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzNEREQzMzNERERERERERERERERERERERERERERERERERERVVVVVVVVERERVVVVVVVVERERVVVVERERERERERERERERVVVVVVVVERERVVVVVVVVVVVVmZmZmZmZmZmZ3d3eIiIiIiIiIiIh3d3dmZmZVVVV3d3eIiIiIiIiZmZmqqqqZmZmqqqqqqqqqqqq7u7vMzMzd3d3u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d7u7u3d3d7u7u3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3dzMzMu7u7qqqqqqqqu7u7zMzMzMzMzMzMzMzMzMzMu7u7zMzMzMzMzMzM3d3dzMzM3d3dzMzMzMzM3d3d3d3d3d3dzMzM3d3d3d3dzMzMzMzMzMzMu7u7u7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqmZmZqqqqmZmZmZmZqqqqmZmZiIiIiIiId3d3d3d3ZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVZmZmd3d3ZmZmZmZmd3d3d3d3ZmZmVVVVVVVVZmZmZmZmd3d3ZmZmd3d3d3d3iIiId3d3iIiIiIiIiIiIiIiId3d3iIiIiIiIqqqqqqqqzMzM3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7uu7u7qqqqu7u7zMzM3d3d3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7uzMzMzMzMu7u7u7u7qqqqqqqqqqqqmZmZmZmZiIiIiIiId3d3iIiIiIiId3d3iIiIiIiImZmZmZmZmZmZmZmZqqqqu7u7u7u7qqqqu7u7qqqqmZmZmZmZmZmZiIiId3d3iIiIVVVVREREREREMzMzMzMzREREREREMzMzREREREREREREREREREREREREREREREREVVVVVVVVREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREVVVVREREREREREREREREREREREREVVVVREREVVVVREREVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVZmZmZmZmiIiId3d3ZmZmZmZmd3d3d3d3iIiIiIiIiIiId3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVMzMzREREVVVVREREVVVVVVVVVVVVREREREREVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVREREREREVVVVVVVVVVVVVVVVREREREREVVVVREREVVVVREREVVVVREREVVVVREREREREREREREREREREREREMzMzMzMzREREREREREREMzMzREREMzMzREREREREREREREREREREREREREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVREREREREVVVVREREVVVVVVVVVVVVREREVVVVVVVVVVVVREREVVVVVVVVVVVVREREREREREREZmZmZmZmVVVVREREREREMzMzMzMzMzMzMzMzMzMzREREREREREREREREVVVVREREREREMzMzMzMzREREZmZmVVVVVVVVVVVVMzMzMzMzREREREREREREREREMzMzREREREREREREREREMzMzREREMzMzREREREREREREREREMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVVVVVVVVVMzMzMzMzREREMzMzMzMzMzMzREREMzMzREREMzMzMzMzREREMzMzMzMzIiIiIiIiIiIiMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzIiIiIiIiMzMzMzMzMzMzREREREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzREREREREREREREREMzMzIiIiMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiMzMzMzMzMzMzREREMzMzMzMzMzMzVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVREREREREREREREREVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmVVVVZmZmVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVZmZmVVVVVVVVZmZmVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3d3d3ZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3ZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3ZmZmd3d3iIiIiIiIiIiId3d3d3d3d3d3d3d3ZmZmZmZmd3d3d3d3d3d3mZmZiIiImZmZiIiImZmZmZmZmZmZiIiIiIiIZmZmVVVVVVVVd3d3VVVVREREVVVVREREVVVVREREVVVVVVVVVVVVREREREREREREREREREREVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVVVVVREREREREREREMzMzMzMzIiIiIiIiMzMzIiIiMzMzMzMzMzMzREREd3d3mZmZqqqqqqqqqqqqmZmZmZmZiIiId3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmVVVVZmZmZmZmZmZmVVVVVVVVREREREREVVVVREREVVVVVVVVVVVVREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVREREVVVVREREVVVVREREVVVVVVVVZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmVVVVZmZmVVVVVVVVREREMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzREREREREREREREREMzMzMzMzMzMzREREREREREREREREREREVVVVREREREREREREREREREREREREVVVVREREVVVVREREVVVVVVVVREREVVVVREREREREVVVVVVVVVVVVVVVVZmZmVVVVd3d3d3d3iIiIiIiIiIiId3d3d3d3ZmZmd3d3iIiImZmZmZmZmZmZqqqqqqqqu7u7u7u7zMzM3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7t3d3d3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3e7u7u7u7u7u7v///+7u7v///////////////+7u7u7u7u7u7u7u7t3d3czMzMzMzLu7u7u7u7u7u8zMzN3d3d3d3d3d3e7u7t3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzN3d3czMzMzMzN3d3czMzMzMzN3d3d3d3czMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u8zMzLu7u6qqqru7u6qqqru7u6qqqqqqqqqqqpmZmZmZmYiIiHd3d2ZmZmZmZmZmZlVVVVVVVWZmZlVVVVVVVWZmZlVVVWZmZmZmZnd3d3d3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d2ZmZmZmZlVVVVVVVWZmZlVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d2ZmZnd3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d4iIiIiIiIiIiJmZmZmZmZmZmZmZmaqqqru7u8zMzO7u7u7u7v///////////////////////////////////////////////////////////////////+7u7v///////////////+7u7v///////////////////////////////////////+7u7v///+7u7u7u7u7u7u7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3e7u7t3d3e7u7u7u7u7u7t3d3e7u7u7u7t3d3d3d3d3d3czMzKqqqqqqqoiIiHd3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d4iIiJmZmZmZmaqqqru7u7u7u7u7u7u7u7u7u6oA//8AAKqqqqqqqqqqqqqqqqqqqqqqqqqqmZmZiIiId3d3d3d3ZmZmREREREREMzMzMzMzREREMzMzMzMzMzMzREREREREREREREREREREREREREREVVVVREREREREMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVREREVVVVREREVVVVREREREREVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmd3d3iIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmVVVVREREVVVVVVVVVVVVZmZmZmZmVVVVREREREREVVVVVVVVREREVVVVREREVVVVVVVVZmZmZmZmd3d3ZmZmZmZmVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmVVVVREREREREVVVVVVVVZmZmVVVVREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVREREVVVVREREMzMzREREMzMzREREREREREREMzMzMzMzREREREREMzMzREREREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVREREVVVVVVVVREREREREVVVVVVVVVVVVVVVVVVVVREREREREREREREREVVVVREREREREREREREREVVVVZmZmZmZmREREMzMzMzMzMzMzMzMzREREREREMzMzREREREREREREREREREREREREMzMzMzMzMzMzZmZmZmZmVVVVVVVVREREMzMzREREREREREREMzMzREREREREMzMzREREREREREREMzMzMzMzREREREREVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzREREVVVVVVVVREREMzMzMzMzMzMzREREMzMzREREMzMzREREREREMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzIiIiMzMzIiIiMzMzMzMzIiIiMzMzIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzREREREREMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiMzMzMzMzMzMzIiIiMzMzREREREREMzMzREREVVVVREREREREMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREZmZmd3d3ZmZmVVVVVVVVVVVVREREVVVVVVVVREREMzMzREREREREVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmVVVVREREREREREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmVVVVVVVVVVVVZmZmVVVVVVVVZmZmVVVVVVVVZmZmVVVVZmZmVVVVVVVVZmZmZmZmVVVVZmZmVVVVZmZmVVVVZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmVVVVZmZmVVVVZmZmVVVVZmZmVVVVZmZmVVVVZmZmZmZmVVVVVVVVZmZmZmZmVVVVVVVVREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3iIiIiIiIiIiIiIiId3d3iIiId3d3ZmZmZmZmd3d3ZmZmZmZmd3d3d3d3d3d3iIiIiIiImZmZmZmZqqqqqqqqmZmZiIiId3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREMzMzVVVVVVVVVVVVREREREREREREVVVVREREVVVVVVVVVVVVREREREREMzMzREREMzMzREREMzMzMzMzMzMzIiIiMzMzIiIiMzMzREREREREREREZmZmmZmZqqqqqqqqqqqqmZmZmZmZiIiId3d3iIiId3d3d3d3ZmZmZmZmVVVVZmZmZmZmZmZmVVVVVVVVZmZmVVVVVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmd3d3iIiId3d3d3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVMzMzREREMzMzREREREREREREMzMzMzMzREREREREREREREREMzMzREREMzMzVVVVVVVVREREMzMzREREREREMzMzREREREREREREREREVVVVVVVVREREREREREREVVVVVVVVREREVVVVREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmd3d3d3d3iIiImZmZmZmZd3d3d3d3d3d3d3d3d3d3mZmZqqqqqqqqu7u7u7u7zMzMzMzMzMzM7u7u7u7u////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7v///////////////////////////////////////////////+7u7t3d3czMzLu7u6qqqqqqqqqqqszMzMzMzN3d3d3d3d3d3d3d3d3d3czMzLu7u7u7u8zMzMzMzLu7u8zMzMzMzMzMzN3d3czMzMzMzLu7u8zMzLu7u8zMzLu7u8zMzLu7u8zMzLu7u8zMzMzMzLu7u7u7u7u7u7u7u8zMzLu7u7u7u8zMzLu7u7u7u6qqqqqqqpmZmaqqqqqqqqqqqpmZmYiIiHd3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiJmZmYiIiIiIiIiIiIiIiJmZmYiIiJmZmYiIiHd3d3d3d3d3d3d3d2ZmZlVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZnd3d2ZmZmZmZmZmZmZmZnd3d3d3d3d3d2ZmZmZmZmZmZnd3d2ZmZmZmZmZmZnd3d4iIiJmZmaqqqqqqqru7u7u7u7u7u93d3e7u7v///////////////////////////////////////////////////+7u7v///////////+7u7v///////////////////////////////////////////////////////////////////////+7u7v///////+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzLu7u7u7u6qqqoiIiHd3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiJmZmaqqqru7u7u7u6qqqqqqqqqqqpmZmZmZmZmZmYiIiJmZmYiIiIiIiJmZmZmZmZmZmbu7u5mZmYiIiHd3d3d3d2ZmZlVVVURERDMzM0RERERERDMzMzMzMzMzMzMzM0RERDMzMzMzM0RERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVURERFVVVVVVVWZmZlVVVVVVVVVVVVVVVWZmZnd3d2ZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVURERERERFVVVURERFVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZoiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d2ZmZmZmZlVVVVVVVVVVVWZmZmZmZlVVVURERERERERERFVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVWZmZmZmZlVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZnd3d2ZmZmZmZnd3d2ZmZlVVVURERERERERERERERFVVVWZmZlVVVVVVVURERERERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERDMzM0RERERERFVVVURERDMzMzMzMzMzMzMzM0RERDMzM0RERERERERERERERERERFVVVVVVVVVVVVVVVVVVVURERFVVVWZmZmZmZmZmZlVVVURERERERERERFVVVURERFVVVVVVVURERFVVVURERFVVVURERFVVVURERERERERERERERERERERERFVVVWZmZmZmZkRERERERDMzM0RERERERDMzM0RERERERERERERERFVVVURERERERERERDMzMzMzM0RERFVVVWZmZmZmZkRERERERERERERERERERERERERERERERDMzM0RERERERERERERERDMzMzMzMzMzM0RERFVVVURERDMzMzMzM0RERDMzMzMzM0RERERERDMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzM0RERERERFVVVVVVVURERDMzM0RERDMzMzMzM0RERDMzM0RERERERDMzM0RERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERERERCIiIjMzMyIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIjMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMyIiIjMzMzMzM0RERERERDMzMzMzM0RERERERERERERERDMzMzMzMzMzMyIiIjMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVWZmZkRERERERDMzM0RERDMzMzMzMzMzMzMzM1VVVVVVVWZmZlVVVWZmZmZmZlVVVWZmZlVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVURERFVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERERERERERFVVVVVVVURERERERDMzMzMzMzMzMzMzMzMzM0RERFVVVWZmZmZmZlVVVVVVVVVVVURERFVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d4iIiIiIiIiIiHd3d3d3d2ZmZmZmZmZmZnd3d3d3d2ZmZmZmZnd3d3d3d4iIiIiIiHd3d3d3d4iIiHd3d4iIiIiIiIiIiIiIiIiIiHd3d3d3d4iIiHd3d3d3d3d3d3d3d2ZmZmZmZnd3d3d3d3d3d4iIiJmZmaqqqqqqqqqqqpmZmZmZmXd3d2ZmZmZmZlVVVVVVVURERGZmZmZmZkRERERERERERERERERERERERERERFVVVVVVVURERERERDMzM0RERERERFVVVVVVVVVVVVVVVURERDMzMzMzM0RERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERHd3d5mZmaqqqqqqqpmZmZmZmYiIiIiIiIiIiIiIiHd3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVURERFVVVWZmZmZmZkRERERERFVVVVVVVWZmZlVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZnd3d4iIiIiIiIiIiHd3d2ZmZnd3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM0RERERERERERFVVVVVVVURERERERERERDMzM0RERERERERERERERERERFVVVURERERERERERFVVVVVVVURERERERFVVVVVVVURERERERFVVVVVVVVVVVWZmZmZmZnd3d4iIiIiIiIiIiJmZmYiIiIiIiHd3d4iIiIiIiJmZmZmZmaqqqru7u8zMzN3d3d3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7d3d3d3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d27u7u7u7vMzMzMzMzMzMy7u7vMzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7vMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMy7u7vMzMy7u7u7u7vMzMy7u7uqqqq7u7uqqqqqqqqqqqq7u7u7u7uqqqqZmZmIiIh3d3eIiIh3d3eIiIiZmZmIiIiZmZmZmZmZmZmZmZmZmZmZmZmIiIiIiIiIiIiIiIiZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmIiIh3d3d3d3d3d3eIiIhmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3eIiIiIiIh3d3d3d3dmZmZVVVVmZmZmZmZ3d3d3d3d3d3eZmZm7u7vMzMzMzMzu7u7d3d3u7u7////u7u7////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////u7u7////////u7u7////u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMy7u7u7u7uqqqqqqqq7u7uqqqqqqqq7u7u7u7uqqqq7u7uqqqqZmZmIiIiZmZmZmZmZmZmZmZmZmZmIiIiIiIiIiIiIiIiIiIiZmZmqqqqqqqq7u7u7u7u7u7u7u7uqqqqZmZlmZmZVVVVVVVVVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzNERERERERERERVVVVVVVVVVVVERERERERVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVERERERERVVVVERERVVVVERERVVVVVVVVVVVVERERVVVVVVVVVVVVmZmZmZmZVVVVmZmZ3d3dmZmZmZmZ3d3d3d3eIiIiIiIiIiIh3d3d3d3dmZmZmZmZmZmZVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERmZmZ3d3dVVVVERERVVVVVVVVmZmZVVVVmZmZVVVVVVVVmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZ3d3dmZmZVVVVVVVVERERVVVVVVVVVVVVmZmZVVVVVVVVVVVVERERERERVVVVERERVVVVERERVVVVVVVVmZmZVVVVVVVVVVVVEREQzMzNERERERERVVVVEREQzMzMzMzNERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVERERVVVVVVVVmZmZmZmZERERVVVVERERVVVVVVVVERERVVVVERERVVVVERERVVVVERERVVVVERERVVVVERERERERERERERERVVVVVVVVVVVVmZmZEREREREREREQzMzMzMzNEREQzMzNERERERERERERERERVVVVERERVVVUzMzMzMzNERERVVVVmZmZmZmZVVVUzMzNERERERERERERVVVVEREREREREREREREREREREREREREREREQzMzMzMzNEREREREREREQzMzMzMzMzMzNEREQzMzNEREQzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzNERERERERVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNEREQzMzNEREREREQzMzMiIiIzMzMzMzMiIiJEREREREQzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREREREQzMzMiIiIzMzMzMzMiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzNERERVVVVEREREREQzMzMzMzMiIiIzMzMzMzMiIiJERERVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVERERVVVVERERERERERERERERVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVEREREREQzMzMzMzNEREREREQzMzMzMzMzMzNERERERERVVVVVVVVERERVVVV3d3d3d3dmZmZVVVVVVVVERERVVVVERERERERVVVV3d3d3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZ3d3dmZmZ3d3dmZmZ3d3d3d3dmZmZ3d3d3d3d3d3d3d3eIiIh3d3eIiIh3d3d3d3d3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3eIiIiIiIiZmZmIiIiIiIiIiIiIiIh3d3eIiIiIiIiIiIiIiIh3d3eZmZmZmZmZmZmqqqq7u7uqqqqZmZmIiIiIiIh3d3dmZmZVVVVVVVVVVVVmZmZVVVVERERERERERERERERERERERERmZmZVVVVEREQzMzNERERERERERERERERVVVVmZmZVVVVEREREREREREREREQzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVEREQzMzNERESIiIiqqqqqqqqqqqqqqqqZmZmIiIiIiIiIiIiIiIh3d3d3d3d3d3dmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZVVVVERERVVVVmZmZERERERERVVVVVVVVVVVVmZmZVVVVmZmZmZmZVVVVVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIh3d3dmZmZmZmZmZmZVVVVmZmZmZmZVVVVVVVVVVVVVVVVEREREREQzMzMzMzMzMzMzMzMzMzNEREQzMzNEREQzMzMzMzNEREQzMzNERERVVVVVVVVVVVVVVVVEREQzMzNERERVVVVERERVVVVERERVVVVERERVVVVVVVVVVVVVVVVERERERERERERERERVVVVVVVVVVVVmZmZmZmZ3d3d3d3eZmZmZmZmZmZmZmZmIiIiIiIh3d3eIiIiIiIiZmZmqqqq7u7vMzMzd3d3d3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u7u7u7u7u3d3d3d3d7u7u3d3d3d3dzMzMzMzM3d3dzMzMzMzMzMzMzMzMzMzMu7u7zMzMzMzMzMzMzMzMzMzM3d3d3d3du7u7u7u7u7u7qqqqqqqqqqqqqqqqu7u7u7u7u7u7u7u7u7u7u7u7zMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7zMzMu7u7u7u7qqqqu7u7u7u7qqqqu7u7u7u7u7u7u7u7u7u7u7u7u7u7zMzMu7u7qqqqmZmZqqqqmZmZmZmZqqqqqqqqqqqqmZmZqqqqqqqqmZmZmZmZqqqqmZmZmZmZmZmZmZmZqqqqqqqqqqqqqqqqmZmZqqqqmZmZmZmZmZmZiIiIiIiId3d3iIiId3d3d3d3d3d3d3d3ZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiId3d3ZmZmZmZmZmZmd3d3d3d3mZmZmZmZqqqqzMzM3d3d7u7u7u7u////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////7u7u////7u7u7u7u////7u7u////7u7u7u7u7u7u7u7u7u7u3d3d3d3dzMzMzMzMu7u7u7u7u7u7zMzMzMzMzMzMu7u7zMzMzMzMu7u7u7u7zMzMu7u7u7u7qqqqmZmZmZmZiIiIiIiId3d3d3d3ZmZmiIiIiIiImZmZiIiImZmZmZmZqqqqqqqqu7u7u7u7zMzMzMzMzMzMzMzMu7u7mZmZd3d3VVVVVVVVREREREREMzMzMzMzMzMzREREREREREREMzMzIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREREREREREREREVVVVVVVVREREREREREREREREREREREREREREREREVVVVVVVVVVVVZmZmVVVVREREREREVVVVREREVVVVVVVVVVVVREREREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmd3d3VVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVREREREREREREZmZmZmZmREREREREMzMzMzMzMzMzMzMzREREREREREREREREREREVVVVVVVVREREVVVVZmZmVVVVVVVVREREVVVVVVVVZmZmVVVVVVVVREREVVVVREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREREREVVVVREREVVVVVVVVZmZmVVVVREREREREREREMzMzREREREREREREREREVVVVREREREREVVVVVVVVREREMzMzMzMzVVVVd3d3ZmZmVVVVREREREREREREREREREREREREREREREREREREREREREREREREREREREREMzMzMzMzVVVVREREMzMzMzMzMzMzMzMzREREREREREREREREREREREREMzMzREREREREMzMzREREMzMzIiIiIiIiIiIiMzMzMzMzREREREREVVVVREREREREMzMzMzMzREREMzMzMzMzMzMzREREMzMzMzMzREREMzMzMzMzMzMzIiIiIiIiMzMzMzMzVVVVMzMzMzMzMzMzMzMzIiIiIiIiMzMzIiIiIiIiMzMzMzMzIiIiMzMzIiIiMzMzIiIiIiIiMzMzREREREREREREREREMzMzMzMzIiIiMzMzMzMzIiIiMzMzMzMzIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzMzMzMzMzIiIiIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREREREMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiMzMzVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVREREVVVVVVVVREREREREREREREREVVVVREREREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmVVVVZmZmVVVVZmZmVVVVZmZmZmZmZmZmd3d3ZmZmVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVREREREREREREREREREREREREVVVVREREVVVVVVVVZmZmZmZmZmZmd3d3ZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmd3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3iIiIiIiId3d3d3d3d3d3ZmZmZmZmZmZmZmZmd3d3d3d3iIiIqqqqqqqqqqqqqqqqmZmZmZmZiIiIiIiIiIiImZmZiIiIiIiImZmZmZmZmZmZqqqqqqqqqqqqmZmZmZmZmZmZiIiId3d3d3d3ZmZmVVVVVVVVZmZmREREREREMzMzMzMzREREVVVVZmZmREREREREMzMzREREREREREREREREVVVVVVVVZmZmREREREREREREREREREREREREREREREREREREREREREREMzMzMzMzREREMzMzREREVVVVREREMzMzMzMzVVVVd3d3mZmZqqqqqqqqmZmZmZmZmZmZmZmZiIiIiIiImZmZiIiIiIiId3d3ZmZmZmZmZmZmd3d3ZmZmZmZmVVVVREREVVVVREREREREREREREREREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmZmZmZmZmZmZmd3d3ZmZmVVVVVVVVVVVVVVVVVVVVREREREREREREREREMzMzREREMzMzREREREREMzMzMzMzREREREREREREREREREREVVVVVVVVREREREREREREREREREREREREREREREREREREVVVVREREREREREREVVVVREREVVVVVVVVVVVVVVVVd3d3d3d3d3d3mZmZmZmZmZmZmZmZiIiId3d3iIiImZmZqqqqqqqqzMzMzMzM7u7u7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////+7u7v///+7u7u7u7u7u7t3d3d3d3czMzN3d3czMzN3d3czMzN3d3d3d3czMzMzMzMzMzLu7u8zMzLu7u8zMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzN3d3czMzKqqqqqqqpmZmZmZmaqqqqqqqqqqqru7u8zMzMzMzMzMzLu7u7u7u7u7u7u7u7u7u8zMzMzMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u8zMzMzMzLu7u7u7u7u7u7u7u7u7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqru7u7u7u6qqqqqqqru7u7u7u7u7u7u7u7u7u6qqqpmZmZmZmYiIiIiIiJmZmYiIiJmZmYiIiHd3d4iIiIiIiIiIiJmZmZmZmZmZmZmZmYiIiIiIiHd3d3d3d3d3d3d3d5mZmZmZmbu7u8zMzMzMzN3d3e7u7u7u7v///////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3czMzLu7u7u7u7u7u7u7u8zMzMzMzMzMzMzMzN3d3czMzMzMzMzMzKqqqqqqqpmZmZmZmXd3d2ZmZlVVVWZmZmZmZnd3d3d3d3d3d3d3d4iIiKqqqqqqqqqqqru7u7u7u8zMzMzMzMzMzKqqqqqqqoiIiHd3d2ZmZlVVVURERDMzMyIiIjMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERFVVVVVVVVVVVURERFVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERFVVVURERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERFVVVURERERERERERERERERERERERFVVVVVVVVVVVWZmZlVVVVVVVXd3d3d3d3d3d3d3d4iIiHd3d4iIiJmZmZmZmXd3d2ZmZnd3d2ZmZmZmZlVVVVVVVVVVVVVVVWZmZlVVVURERERERFVVVVVVVVVVVWZmZnd3d3d3d2ZmZlVVVVVVVWZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZmZmZnd3d2ZmZlVVVURERFVVVVVVVURERFVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d2ZmZlVVVURERERERDMzM0RERERERERERERERERERERERERERFVVVVVVVVVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVWZmZlVVVURERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVURERERERFVVVXd3d2ZmZkRERERERERERERERERERERERFVVVURERFVVVVVVVVVVVVVVVVVVVURERERERDMzM1VVVXd3d2ZmZkRERERERDMzM0RERFVVVURERFVVVURERERERFVVVURERFVVVURERERERERERERERERERERERFVVVTMzM0RERDMzM0RERDMzMzMzM0RERERERERERDMzM0RERDMzM0RERERERERERDMzMyIiIiIiIiIiIjMzMzMzM0RERERERFVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzM0RERERERDMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzM0RERERERERERDMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMyIiIjMzMzMzM0RERERERERERDMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMyIiIjMzMyIiIiIiIjMzMyIiIjMzMzMzM0RERERERERERERERERERERERFVVVURERFVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERFVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZnd3d2ZmZnd3d2ZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZnd3d2ZmZmZmZmZmZnd3d2ZmZnd3d3d3d2ZmZnd3d3d3d3d3d3d3d2ZmZmZmZnd3d3d3d2ZmZnd3d2ZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZnd3d2ZmZnd3d3d3d3d3d3d3d4iIiIiIiIiIiHd3d3d3d3d3d3d3d2ZmZnd3d2ZmZmZmZnd3d3d3d4iIiIiIiIiIiJmZmZmZmZmZmZmZmaqqqpmZmZmZmZmZmaqqqpmZmZmZmZmZmZmZmaqqqqqqqpmZmZmZmZmZmZmZmZmZmYiIiIiIiHd3d3d3d2ZmZmZmZmZmZmZmZkRERERERDMzM0RERFVVVURERFVVVWZmZkRERERERERERERERERERERERFVVVURERGZmZmZmZkRERERERERERERERERERERERERERERERERERERERERERERERERERERERERERFVVVVVVVURERDMzMzMzM0RERERERGZmZoiIiJmZmZmZmZmZmYiIiIiIiIiIiJmZmZmZmYiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d3d3d2ZmZlVVVVVVVURERERERERERERERERERERERFVVVVVVVVVVVWZmZnd3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d2ZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVURERFVVVVVVVURERDMzM0RERERERERERERERERERERERDMzM0RERDMzM0RERERERERERERERFVVVVVVVVVVVURERERERERERFVVVURERERERFVVVURERERERFVVVVVVVURERGZmZmZmZmZmZnd3d3d3d4iIiJmZmZmZmZmZmZmZmZmZmZmZmZmZmaqqqszMzN3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3MzMzd3d3MzMzMzMzMzMy7u7vMzMy7u7u7u7vMzMzMzMy7u7uqqqqqqqqqqqq7u7u7u7vMzMy7u7vMzMy7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7uqqqqqqqq7u7u7u7u7u7u7u7vMzMy7u7u7u7u7u7u7u7vMzMy7u7vMzMy7u7vMzMy7u7vMzMzMzMy7u7vMzMy7u7u7u7uqqqq7u7uqqqqqqqqqqqq7u7u7u7u7u7u7u7u7u7u7u7u7u7uqqqqqqqq7u7u7u7u7u7vMzMzMzMy7u7u7u7uqqqqqqqqqqqqZmZmqqqq7u7uqqqqqqqqZmZmZmZmZmZmZmZmZmZmqqqqZmZmZmZmIiIiIiIh3d3eIiIiZmZmqqqq7u7vd3d3u7u7u7u7////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7u7u7u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3MzMy7u7u7u7u7u7u7u7vMzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7uqqqqIiIiIiIiIiIh3d3d3d3dmZmZmZmZ3d3d3d3eIiIiZmZmqqqqqqqq7u7u7u7u7u7u7u7u7u7vMzMzMzMy7u7uZmZlmZmZVVVVEREQzMzMiIiIiIiIzMzMiIiIzMzMiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMiIiIiIiIzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzNERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVEREQzMzNVVVVEREQzMzMzMzMzMzMzMzMzMzNEREQzMzNERERERERERERERERERERERERVVVVERERERERERERVVVVERERVVVVVVVVERERVVVVEREREREREREQzMzNERERERERERERERERERERERERVVVVERERVVVVERERERERVVVVVVVVVVVV3d3d3d3d3d3d3d3eIiIh3d3d3d3eIiIiZmZmZmZmIiIh3d3eIiIh3d3dmZmZ3d3d3d3dmZmZVVVVVVVVVVVVVVVVERERERERVVVVVVVVmZmaIiIiIiIh3d3dmZmZmZmZVVVVmZmZVVVVmZmZ3d3dmZmZmZmZ3d3d3d3d3d3dmZmZERERVVVVERERERERVVVVVVVVVVVVERERERERVVVVERERERERVVVVERERVVVVVVVVVVVVmZmZmZmZVVVVERERVVVVERERVVVVERERERERERERERERERERERERERERVVVVVVVVVVVVmZmZVVVVmZmZVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERVVVVVVVVmZmZmZmZVVVVVVVVVVVVERERmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZVVVVERERERERERERVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVUzMzNERERVVVV3d3dmZmZVVVVERERERERERERERERVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVERERERERERERERERVVVVEREQzMzNEREQzMzNERERERERERERERERERERVVVVEREQzMzNEREQzMzNEREQzMzMiIiIiIiIiIiIzMzMzMzNERERERERVVVVEREQzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIzMzNEREREREQzMzMiIiIzMzMzMzMiIiIiIiIiIiIiIiIzMzMiIiIiIiIzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzNVVVVEREQzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMiIiIiIiIzMzMiIiIzMzMzMzMiIiIzMzMiIiIzMzMzMzNEREQzMzNEREQzMzNERERERERERERVVVVERERERERERERVVVVVVVVERERVVVVmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZ3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZ3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3eIiIiIiIh3d3eIiIh3d3d3d3dmZmZ3d3dmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3eIiIiIiIh3d3d3d3d3d3eIiIiIiIiZmZmqqqqqqqqqqqqqqqqqqqqZmZmZmZmZmZmZmZmIiIh3d3eIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3eIiIh3d3d3d3dmZmZERERERERVVVVVVVVVVVVERERmZmZmZmZVVVVERERERERERERERERVVVVERERVVVVVVVVmZmZVVVVERERVVVVERERERERERERERERERERVVVVmZmZVVVVERERERERERERERERVVVVVVVVEREQzMzNERERERERERERERERmZmZ3d3eIiIiZmZmIiIiIiIiIiIiIiIiZmZmIiIiIiIiIiIiIiIiIiIh3d3eIiIiIiIh3d3d3d3d3d3dmZmZVVVVEREREREREREREREQzMzNVVVVERERVVVVmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIhmZmZmZmZmZmZVVVVmZmZ3d3dmZmZmZmZVVVVmZmZmZmZmZmZVVVVVVVVVVVVERERVVVVEREREREREREREREREREQzMzNERERERERERERERERERERERERVVVVERERERERERERERERVVVVERERVVVVERERVVVVERERVVVVERERVVVVVVVVmZmZmZmZ3d3d3d3d3d3eIiIiIiIiIiIiZmZmqqqqqqqrMzMzMzMzu7u7u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3d3d3d3d3d3d3d3d3d7u7u3d3d3d3d7u7u3d3d3d3d3d3dzMzMzMzMzMzMzMzMu7u7u7u7zMzMzMzM3d3dzMzMzMzMu7u7u7u7u7u7qqqqu7u7u7u7zMzMzMzMzMzMzMzMu7u7u7u7u7u7qqqqu7u7qqqqqqqqqqqqqqqqqqqqu7u7u7u7zMzMzMzMu7u7zMzMzMzMzMzMzMzMzMzM3d3dzMzM3d3dzMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7zMzMu7u7u7u7u7u7u7u7u7u7u7u7qqqqqqqqu7u7u7u7zMzMzMzMzMzMzMzMzMzMu7u7u7u7qqqqu7u7u7u7u7u7u7u7zMzMu7u7qqqqqqqqmZmZmZmZqqqqmZmZmZmZmZmZmZmZmZmZqqqqu7u7zMzM7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////7u7u////////////////////////////7u7u7u7u7u7u7u7u7u7u7u7u////7u7u////7u7u7u7u7u7u3d3dzMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7qqqqqqqqiIiImZmZiIiIiIiId3d3iIiImZmZmZmZqqqqmZmZmZmZqqqqu7u7u7u73d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMu7u7mZmZd3d3REREREREMzMzMzMzMzMzMzMzMzMzREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzREREREREREREREREREREVVVVREREREREVVVVVVVVVVVVZmZmVVVVVVVVREREVVVVREREREREREREREREMzMzREREMzMzMzMzMzMzREREMzMzREREREREREREREREVVVVVVVVREREVVVVREREREREREREREREREREREREREREREREREREMzMzREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREVVVVZmZmd3d3ZmZmZmZmVVVVd3d3iIiImZmZd3d3ZmZmd3d3d3d3mZmZiIiId3d3iIiId3d3d3d3ZmZmREREREREREREREREVVVVREREZmZmd3d3d3d3iIiId3d3d3d3ZmZmZmZmVVVVZmZmZmZmZmZmZmZmd3d3ZmZmZmZmVVVVREREREREREREREREREREREREVVVVVVVVVVVVREREREREVVVVVVVVREREVVVVVVVVVVVVZmZmVVVVVVVVREREREREREREREREREREVVVVVVVVREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVREREZmZmZmZmZmZmZmZmVVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmd3d3ZmZmZmZmVVVVVVVVZmZmZmZmZmZmVVVVVVVVREREVVVVREREREREVVVVVVVVREREVVVVZmZmZmZmVVVVVVVVREREREREZmZmd3d3d3d3VVVVREREVVVVVVVVZmZmVVVVVVVVZmZmVVVVREREVVVVVVVVVVVVREREVVVVREREREREREREVVVVREREREREMzMzREREREREREREREREVVVVREREREREREREREREMzMzREREMzMzMzMzMzMzIiIiIiIiMzMzREREVVVVREREREREVVVVREREMzMzREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiREREREREMzMzMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREREREMzMzIiIiMzMzIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzMzMzREREVVVVMzMzREREZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmVVVVZmZmd3d3d3d3ZmZmd3d3ZmZmd3d3d3d3ZmZmZmZmd3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3ZmZmZmZmZmZmd3d3ZmZmZmZmd3d3d3d3iIiIiIiIiIiId3d3iIiId3d3d3d3d3d3d3d3d3d3iIiIiIiImZmZqqqqmZmZmZmZmZmZqqqqmZmZmZmZd3d3ZmZmVVVVZmZmZmZmZmZmd3d3ZmZmd3d3d3d3iIiImZmZiIiIiIiId3d3ZmZmVVVVVVVVZmZmVVVVREREREREVVVVZmZmVVVVVVVVREREVVVVREREVVVVREREVVVVZmZmZmZmZmZmREREREREVVVVREREVVVVREREVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREMzMzREREREREREREREREREREZmZmd3d3iIiImZmZmZmZmZmZiIiIiIiImZmZiIiIiIiIiIiIiIiId3d3iIiIiIiIiIiIiIiIZmZmZmZmVVVVVVVVVVVVREREREREVVVVVVVVREREZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3iIiId3d3iIiIZmZmZmZmVVVVZmZmZmZmZmZmZmZmd3d3ZmZmZmZmd3d3ZmZmZmZmVVVVVVVVREREREREVVVVREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVREREZmZmZmZmZmZmZmZmZmZmd3d3iIiIiIiIiIiId3d3iIiImZmZqqqqzMzM3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7t3d3d3d3d3d3d3d3d3d3e7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3d3d3d3d3e7u7u7u7t3d3e7u7t3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzN3d3d3d3czMzLu7u7u7u7u7u7u7u8zMzMzMzMzMzLu7u7u7u7u7u7u7u6qqqqqqqqqqqru7u7u7u7u7u6qqqqqqqqqqqqqqqru7u7u7u7u7u8zMzMzMzLu7u8zMzMzMzMzMzN3d3czMzN3d3czMzMzMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u8zMzLu7u7u7u7u7u6qqqru7u6qqqqqqqru7u7u7u8zMzMzMzLu7u8zMzMzMzLu7u8zMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u6qqqqqqqpmZmZmZmaqqqqqqqru7u8zMzMzMzO7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7v///////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7u7u7u7u7u7u7v///+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7u7u7szMzMzMzMzMzMzMzMzMzMzMzLu7u6qqqqqqqqqqqqqqqpmZmYiIiHd3d3d3d3d3d5mZmZmZmbu7u7u7u7u7u7u7u8zMzMzMzN3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzLu7u6qqqoiIiGZmZmZmZlVVVURERFVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZlVVVURERFVVVVVVVURERDMzM0RERDMzM0RERERERDMzM0RERERERERERERERERERDMzM1VVVURERFVVVURERERERFVVVURERFVVVURERERERERERERERERERDMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERERERERERERERERERFVVVVVVVVVVVVVVVURERERERERERERERERERDMzM0RERERERERERERERERERERERERERERERERERERERERERDMzMzMzMzMzM0RERDMzMzMzM0RERERERERERFVVVVVVVWZmZlVVVVVVVXd3d5mZmXd3d1VVVVVVVXd3d3d3d4iIiHd3d3d3d4iIiHd3d4iIiGZmZlVVVURERERERERERDMzM0RERFVVVWZmZnd3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZkRERERERERERERERERERDMzM0RERFVVVURERFVVVVVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVURERERERERERDMzM0RERERERFVVVURERFVVVURERERERERERFVVVVVVVWZmZmZmZlVVVWZmZmZmZmZmZmZmZlVVVURERGZmZmZmZmZmZmZmZlVVVVVVVVVVVURERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZlVVVURERFVVVURERFVVVURERFVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVURERGZmZoiIiGZmZkRERERERFVVVURERFVVVVVVVVVVVURERFVVVWZmZlVVVVVVVURERERERERERFVVVURERERERFVVVURERERERERERFVVVVVVVURERERERERERFVVVURERERERERERDMzMzMzMzMzMzMzMzMzMyIiIiIiIkRERERERERERERERERERFVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzM0RERERERDMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMyIiIiIiIjMzMyIiIjMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIiIiIjMzM0RERERERERERCIiIjMzMyIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzM0RERERERDMzMzMzMyIiIjMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzM0RERFVVVURERERERGZmZlVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVWZmZlVVVVVVVWZmZlVVVURERGZmZmZmZmZmZnd3d4iIiHd3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVURERFVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVURERFVVVURERERERFVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVWZmZlVVVWZmZlVVVWZmZmZmZnd3d3d3d2ZmZnd3d2ZmZnd3d2ZmZnd3d3d3d3d3d2ZmZmZmZnd3d3d3d2ZmZnd3d3d3d3d3d3d3d4iIiHd3d3d3d4iIiHd3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiJmZmZmZmZmZmZmZmYiIiIiIiIiIiHd3d1VVVVVVVURERFVVVXd3d2ZmZnd3d2ZmZnd3d3d3d4iIiHd3d4iIiHd3d2ZmZnd3d2ZmZmZmZnd3d1VVVURERDMzM0RERFVVVWZmZmZmZlVVVURERFVVVVVVVVVVVVVVVVVVVWZmZnd3d2ZmZmZmZlVVVURERERERERERFVVVVVVVVVVVVVVVVVVVURERFVVVVVVVWZmZlVVVWZmZlVVVVVVVURERDMzM0RERERERERERERERERERERERGZmZoiIiJmZmYiIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZnd3d2ZmZmZmZmZmZmZmZnd3d3d3d4iIiHd3d4iIiHd3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVURERFVVVVVVVVVVVVVVVURERERERDMzM0RERERERFVVVURERERERDMzM0RERERERERERERERFVVVVVVVURERFVVVWZmZlVVVWZmZmZmZmZmZnd3d3d3d4iIiIiIiJmZmaqqqru7u7u7u6qqqqqqqszMzN3d3f///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMzMzMzMzMzd3d3d3d3d3d3MzMzMzMzMzMzMzMzMzMzMzMzd3d3d3d3MzMzMzMzMzMzMzMy7u7u7u7uqqqqqqqqqqqqqqqq7u7u7u7vMzMy7u7uqqqq7u7u7u7u7u7vMzMzMzMy7u7u7u7vMzMzMzMzMzMy7u7vMzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7uqqqqqqqqqqqqqqqq7u7u7u7vMzMzMzMzMzMzd3d3MzMzMzMzMzMzMzMy7u7u7u7uqqqqqqqqZmZmqqqqZmZm7u7u7u7vMzMzu7u7u7u7////////////////////////////////////////////////////////u7u7////////////////////////////////////////u7u7////u7u7u7u7////u7u7MzMzd3d3u7u7u7u7////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMy7u7u7u7uqqqqqqqqZmZmZmZmIiIiZmZmIiIiIiIh3d3d3d3eIiIiZmZmZmZmZmZmZmZmqqqqqqqq7u7u7u7u7u7vMzMzMzMy7u7u7u7uqqqqqqqqZmZmZmZl3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZVVVVmZmZmZmZVVVVmZmZ3d3dmZmZmZmZmZmZVVVVVVVVmZmZVVVVVVVVVVVVEREREREREREREREREREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzNERERVVVVVVVVVVVVEREREREREREREREREREQzMzNEREREREREREREREQzMzNEREREREREREQzMzNEREQzMzMzMzNEREQzMzNEREREREREREQzMzNERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVmZmZmZmZ3d3d3d3eIiIhmZmZ3d3d3d3d3d3dmZmZVVVVERERERERERERERERVVVVmZmZmZmZ3d3dmZmZ3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3dmZmZERERERERVVVVVVVVEREREREQzMzNERERERERVVVVERERERERVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZ3d3d3d3dmZmZVVVVVVVV3d3d3d3dVVVVERERERERVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZERERERERERERERERERERERERVVVVERERVVVVmZmZVVVVVVVVEREQzMzNERERERERERERVVVVVVVVERERERERVVVVVVVVVVVVERERVVVVVVVVVVVVEREREREREREREREREREQzMzNEREQzMzMiIiIzMzMzMzMzMzNERERVVVVEREQzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzNEREREREREREREREQzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMiIiIzMzMzMzNEREREREREREQzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzNEREREREQzMzMzMzMiIiIzMzMiIiIiIiIzMzMiIiIzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERVVVVERERERERERERERERERERERERVVVVmZmZmZmZVVVVVVVVmZmZmZmZVVVVVVVVmZmZmZmZmZmaIiIh3d3d3d3dmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVVVVVERERERERVVVVERERVVVVERERVVVVERERVVVVERERVVVVVVVVVVVVmZmZVVVVmZmZVVVVVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERERERERERERERVVVVVVVVERERERERVVVVERERVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3d3d3eIiIiIiIiZmZmIiIiZmZmZmZmZmZmZmZmZmZmIiIiIiIh3d3dmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZ3d3d3d3dmZmZ3d3d3d3d3d3d3d3eIiIiIiIh3d3dmZmZmZmZmZmZ3d3d3d3dVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVV3d3dmZmZmZmZVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZmZmZVVVVVVVVEREREREREREQzMzNERERERERmZmZ3d3eIiIiZmZmZmZmZmZmIiIiIiIiIiIiIiIiZmZmIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3dmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIh3d3eIiIh3d3dmZmZ3d3dmZmZ3d3dmZmZVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVERERERERVVVVERERERERERERERERERERERERERERERERERERERERERERERERERERVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3eIiIiIiIiIiIiZmZmqqqqqqqrMzMzMzMzd3d3d3d3d3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u3d3d7u7u3d3d7u7u3d3d7u7u7u7u3d3d7u7u7u7u3d3d7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzMzMzMzMzM3d3d3d3d3d3dzMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3du7u7u7u7qqqqqqqqqqqqqqqqu7u7u7u7qqqqqqqqu7u7zMzMu7u7u7u7u7u7u7u7zMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7zMzMu7u7zMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7qqqqqqqqqqqqqqqqu7u7u7u7u7u7qqqqu7u7qqqqmZmZmZmZmZmZmZmZqqqqu7u7zMzMzMzMzMzM3d3dzMzMzMzMu7u7u7u7qqqqqqqqqqqqmZmZqqqqqqqqu7u73d3d3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////3d3d7u7u7u7u3d3dzMzMzMzM3d3d3d3d7u7u////////////////7u7u////////////////////////////////////////////7u7u7u7u3d3d7u7u3d3d3d3d7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3dzMzMzMzMu7u7u7u7u7u7qqqqqqqqqqqqmZmZqqqqmZmZmZmZmZmZiIiIiIiIiIiId3d3ZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmiIiImZmZqqqqqqqqu7u7u7u7u7u7u7u7qqqqmZmZiIiIiIiImZmZd3d3d3d3d3d3ZmZmVVVVZmZmZmZmVVVVZmZmZmZmZmZmd3d3iIiId3d3d3d3d3d3VVVVZmZmd3d3ZmZmVVVVVVVVVVVVREREREREREREMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVZmZmREREREREREREREREVVVVREREVVVVVVVVZmZmZmZmd3d3ZmZmZmZmZmZmZmZmiIiIiIiId3d3VVVVREREREREVVVVVVVVZmZmZmZmZmZmd3d3ZmZmd3d3d3d3ZmZmZmZmVVVVZmZmZmZmZmZmREREREREVVVVVVVVREREREREREREREREREREVVVVVVVVVVVVVVVVZmZmd3d3d3d3ZmZmZmZmZmZmVVVVREREREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVd3d3ZmZmVVVVREREREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmREREMzMzVVVVREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVd3d3d3d3VVVVVVVVREREVVVVREREREREREREVVVVREREREREVVVVVVVVVVVVREREREREREREREREVVVVREREREREREREREREVVVVREREREREVVVVVVVVVVVVREREVVVVVVVVVVVVREREVVVVREREREREMzMzREREMzMzMzMzREREREREVVVVREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVVVVVREREREREMzMzMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzIiIiMzMzMzMzIiIiIiIiMzMzREREREREREREMzMzMzMzIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzIiIiMzMzMzMzMzMzREREVVVVREREMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREREREMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiMzMzIiIiIiIiMzMzMzMzIiIiMzMzREREMzMzMzMzREREVVVVVVVVMzMzMzMzMzMzMzMzMzMzVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREREREZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREREREREREREREVVVVREREVVVVREREREREMzMzMzMzMzMzMzMzREREREREVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmVVVVZmZmVVVVZmZmVVVVZmZmVVVVVVVVZmZmVVVVZmZmVVVVVVVVZmZmVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmd3d3d3d3d3d3iIiIiIiIiIiId3d3d3d3d3d3ZmZmZmZmd3d3d3d3iIiImZmZmZmZmZmZqqqqqqqqqqqqmZmZiIiId3d3d3d3VVVVREREREREREREREREREREVVVVZmZmZmZmZmZmZmZmd3d3d3d3ZmZmd3d3ZmZmd3d3d3d3mZmZiIiId3d3ZmZmZmZmZmZmZmZmd3d3ZmZmVVVVVVVVZmZmZmZmZmZmVVVVVVVVd3d3iIiIZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmREREVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmiIiIZmZmVVVVVVVVREREREREREREREREREREREREZmZmd3d3d3d3iIiImZmZiIiIiIiIiIiIiIiImZmZmZmZiIiIiIiId3d3iIiIiIiId3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZiIiIiIiIiIiIiIiImZmZmZmZiIiIiIiIiIiIiIiIiIiId3d3iIiId3d3d3d3d3d3ZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVREREVVVVVVVVVVVVVVVVREREREREVVVVREREREREVVVVVVVVREREREREVVVVVVVVZmZmZmZmd3d3d3d3iIiIiIiImZmZmZmZmZmZmZmZqqqqqqqqu7u73d3d7u7u7u7u7u7u////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3czMzN3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzLu7u6qqqpmZmZmZmaqqqqqqqru7u7u7u7u7u8zMzLu7u7u7u8zMzMzMzLu7u7u7u7u7u7u7u8zMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u7u7u6qqqqqqqqqqqqqqqru7u7u7u7u7u7u7u6qqqqqqqqqqqqqqqqqqqqqqqru7u7u7u7u7u7u7u6qqqqqqqpmZmZmZmYiIiJmZmaqqqru7u7u7u8zMzMzMzMzMzLu7u6qqqqqqqpmZmYiIiJmZmZmZmbu7u7u7u8zMzN3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7szMzMzMzO7u7t3d3bu7u6qqqqqqqszMzO7u7v///////////////////////////////////////////////+7u7v///////////+7u7v///+7u7t3d3d3d3d3d3d3d3czMzN3d3d3d3czMzMzMzLu7u7u7u6qqqpmZmaqqqpmZmZmZmZmZmZmZmYiIiHd3d3d3d2ZmZnd3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d3d3d3d3d3d3d5mZmaqqqqqqqqqqqqqqqru7u6qqqqqqqpmZmYiIiIiIiJmZmZmZmXd3d3d3d4iIiHd3d2ZmZmZmZnd3d2ZmZmZmZnd3d2ZmZmZmZnd3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVURERDMzMzMzMzMzMzMzMyIiIiIiIjMzMyIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzM0RERERERDMzM0RERERERFVVVURERFVVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVURERFVVVVVVVURERFVVVVVVVWZmZlVVVWZmZmZmZmZmZnd3d3d3d4iIiJmZmZmZmXd3d2ZmZlVVVVVVVWZmZmZmZmZmZmZmZlVVVWZmZnd3d2ZmZnd3d2ZmZmZmZmZmZkRERERERERERERERFVVVURERERERERERFVVVWZmZlVVVVVVVVVVVWZmZmZmZnd3d3d3d2ZmZmZmZmZmZmZmZjMzM0RERDMzM0RERERERERERFVVVURERFVVVURERFVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZkRERERERFVVVVVVVURERFVVVURERFVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVWZmZmZmZnd3d1VVVVVVVVVVVURERERERERERFVVVWZmZlVVVVVVVURERFVVVVVVVWZmZlVVVWZmZmZmZmZmZoiIiHd3d1VVVVVVVURERFVVVURERFVVVVVVVVVVVURERERERERERERERERERFVVVVVVVURERERERFVVVWZmZmZmZkRERERERDMzM0RERERERFVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVURERERERFVVVVVVVVVVVVVVVVVVVURERERERERERERERERERDMzM0RERFVVVURERERERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERDMzMzMzMyIiIjMzMyIiIjMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERFVVVURERDMzMyIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVVVVVURERDMzMyIiIiIiIjMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMyIiIjMzM0RERFVVVURERERERDMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVURERDMzMzMzMzMzM1VVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZlVVVVVVVURERGZmZnd3d1VVVVVVVURERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERERERDMzM0RERDMzM0RERERERERERERERERERFVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZlVVVWZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVURERFVVVURERERERERERFVVVVVVVVVVVWZmZmZmZnd3d4iIiIiIiIiIiHd3d4iIiHd3d2ZmZnd3d2ZmZlVVVWZmZnd3d3d3d4iIiIiIiJmZmZmZmZmZmZmZmXd3d3d3d2ZmZmZmZlVVVVVVVURERERERERERERERFVVVWZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZnd3d3d3d2ZmZnd3d4iIiHd3d1VVVVVVVVVVVVVVVVVVVWZmZnd3d3d3d2ZmZmZmZlVVVWZmZmZmZmZmZoiIiHd3d1VVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d3d3d2ZmZlVVVWZmZlVVVXd3d4iIiHd3d2ZmZmZmZmZmZlVVVURERERERDMzM0RERFVVVVVVVVVVVVVVVWZmZoiIiIiIiIiIiIiIiJmZmZmZmZmZmYiIiIiIiIiIiIiIiHd3d3d3d4iIiIiIiJmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmaqqqpmZmaqqqpmZmZmZmZmZmZmZmYiIiJmZmYiIiIiIiHd3d3d3d4iIiJmZmYiIiIiIiHd3d3d3d3d3d2ZmZlVVVWZmZmZmZmZmZmZmZlVVVVVVVWZmZnd3d2ZmZmZmZlVVVVVVVWZmZmZmZnd3d3d3d3d3d4iIiIiIiKqqqqqqqqqqqru7u6qqqru7u8zMzMzMzN3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3u7u7d3d3u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3MzMzd3d3d3d3d3d3MzMzd3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMy7u7u7u7u7u7uqqqqqqqqZmZmZmZmqqqq7u7u7u7vMzMzMzMzd3d3MzMzd3d3MzMzMzMzMzMzMzMzMzMy7u7vMzMzMzMzMzMzMzMzMzMzMzMzMzMyqqqq7u7uqqqq7u7u7u7u7u7u7u7u7u7u7u7uqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqq7u7uqqqqqqqqqqqqZmZmZmZmZmZmZmZmqqqqqqqq7u7uqqqqqqqqZmZmZmZmZmZmIiIiZmZmZmZmqqqrMzMzMzMzu7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////d3d2qqqq7u7vd3d3d3d2qqqqZmZmqqqrMzMzu7u7u7u7////////////////////u7u7////////////////////////////////u7u7////d3d27u7uZmZmIiIiZmZmqqqq7u7u7u7vMzMy7u7u7u7u7u7u7u7uqqqqZmZmZmZmZmZmIiIh3d3dmZmZmZmZVVVVmZmZmZmZ3d3dmZmZmZmZmZmZ3d3eIiIiIiIiZmZmZmZmZmZmqqqqqqqqqqqqZmZmqqqqqqqqZmZmZmZmqqqqZmZmqqqqqqqqqqqqIiIiZmZmZmZmZmZmIiIh3d3eZmZmIiIiIiIiIiIh3d3dmZmZVVVVVVVVVVVVERERERERERERERERERERVVVVEREREREQzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzNERERVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVERERERERERERERERVVVVERERVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVERERERERVVVVmZmZVVVVVVVVVVVV3d3dmZmZ3d3eIiIiqqqqZmZmIiIh3d3dVVVVmZmZVVVVmZmZVVVVVVVVmZmZmZmZ3d3d3d3d3d3d3d3dmZmZVVVVEREREREREREREREREREREREREREQzMzNmZmZmZmZVVVVERERERERmZmZmZmZmZmZ3d3dmZmZmZmZmZmZEREQzMzNERERERERERERERERERERERERVVVVVVVVERERERERERERVVVVVVVV3d3d3d3d3d3dmZmZmZmZmZmZVVVVmZmZmZmZmZmZERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVV3d3dmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVERERVVVVVVVVERERERERVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZ3d3d3d3dmZmZERERERERVVVVVVVVERERVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVmZmaIiIh3d3dVVVVVVVVEREREREQzMzNERERERERVVVVmZmZVVVVERERVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVmZmaIiIh3d3dVVVVVVVVERERERERVVVVERERERERERERERERVVVVVVVVVVVVVVVUzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzNVVVVVVVVEREQzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMiIiIiIiIzMzMzMzNEREREREREREQzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVVVVVVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzNERERVVVVERERVVVVVVVVEREREREQzMzMzMzMzMzMiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERVVVVmZmZVVVVERERVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVERERVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZVVVV3d3dmZmZVVVVVVVVVVVVERERERERERERERERVVVVERERVVVVVVVVERERVVVVVVVVERERVVVVVVVVVVVVERERERERVVVVVVVVVVVVERERVVVVERERERERVVVVERERERERERERERERVVVVVVVVmZmZmZmZmZmZVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVERERERERERERERERERERERERVVVVVVVVVVVVmZmZmZmZ3d3d3d3eIiIh3d3d3d3d3d3d3d3dmZmZmZmZmZmZVVVVVVVVmZmZ3d3d3d3eIiIiIiIiIiIiIiIh3d3d3d3dVVVVERERERERERERERERVVVVVVVVVVVVERERERERVVVVmZmZVVVVmZmZmZmZmZmZVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVVVVVmZmZ3d3d3d3d3d3dmZmZVVVVVVVVVVVVmZmaIiIh3d3dmZmZVVVVVVVVVVVVVVVVERERERERVVVVmZmZmZmZmZmZVVVVVVVVmZmZVVVVmZmZVVVVVVVVmZmZ3d3d3d3dVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVERERVVVVmZmZmZmZ3d3eIiIiIiIiZmZmIiIiIiIiZmZmIiIiZmZmIiIiIiIiIiIiIiIiZmZmZmZmqqqqZmZmZmZmZmZmZmZmqqqqZmZmqqqqZmZmqqqqZmZmZmZmqqqqZmZmZmZmIiIiIiIh3d3eIiIiZmZmqqqqqqqqZmZmZmZmIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIh3d3d3d3eIiIiIiIiZmZmIiIiZmZmZmZmqqqqqqqq7u7uqqqqqqqqqqqqqqqq7u7vMzMzd3d3u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////u7u7///////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u3d3d3d3d7u7u3d3d3d3d7u7u7u7u7u7u3d3d7u7u3d3d3d3dzMzMzMzMzMzM3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u73d3du7u7qqqqqqqqqqqqu7u7u7u7u7u7zMzMu7u7zMzM3d3d3d3dzMzM3d3dzMzM3d3dzMzMzMzMzMzMzMzMzMzMzMzM3d3dzMzMu7u7u7u7u7u7u7u7qqqqu7u7u7u7zMzMzMzMu7u7u7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqqqqqmZmZqqqqqqqqqqqqqqqqmZmZqqqqqqqqqqqqqqqqqqqqmZmZmZmZmZmZmZmZmZmZiIiIiIiIiIiImZmZmZmZqqqqu7u7zMzM3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////3d3dqqqqqqqq3d3d7u7uu7u7mZmZzMzM3d3d7u7u////////////////////////////////////////////////////7u7u3d3d3d3dqqqqiIiId3d3d3d3d3d3iIiImZmZqqqqqqqqqqqqu7u7u7u7qqqqmZmZmZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZqqqqu7u7qqqqu7u7u7u7u7u7u7u7u7u7u7u7u7u7qqqqu7u7qqqqqqqqqqqqmZmZmZmZqqqqu7u7qqqqqqqqu7u7qqqqmZmZiIiIiIiIqqqqmZmZmZmZqqqqmZmZiIiId3d3REREREREREREMzMzMzMzREREMzMzREREREREVVVVREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREREREREREREREREREREREMzMzREREREREMzMzMzMzMzMzIiIiREREREREMzMzMzMzMzMzMzMzREREREREREREREREZmZmZmZmd3d3d3d3ZmZmVVVVVVVVREREREREREREREREREREREREREREREREVVVVVVVVREREVVVVVVVVVVVVREREREREREREREREREREREREREREREREVVVVREREVVVVZmZmZmZmd3d3iIiImZmZiIiId3d3d3d3d3d3d3d3ZmZmVVVVZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmREREMzMzREREREREREREREREMzMzREREREREVVVVREREMzMzREREVVVVZmZmd3d3ZmZmd3d3VVVVZmZmVVVVMzMzREREMzMzREREREREREREVVVVREREREREREREREREVVVVVVVVVVVVd3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmVVVVREREREREREREREREVVVVREREVVVVVVVVZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3VVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVZmZmVVVVVVVVZmZmd3d3d3d3iIiIiIiIVVVVREREREREVVVVREREMzMzMzMzREREREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmd3d3d3d3REREREREVVVVVVVVREREREREREREREREREREREREVVVVVVVVVVVVVVVVREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVVVVVREREREREMzMzMzMzIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzVVVVZmZmREREMzMzREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREREREREREREREREREREREREREMzMzMzMzMzMzIiIiMzMzREREREREMzMzREREVVVVZmZmVVVVVVVVREREVVVVREREREREMzMzMzMzMzMzIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREVVVVZmZmZmZmZmZmVVVVVVVVVVVVREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVREREVVVVREREREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmVVVVZmZmd3d3d3d3ZmZmZmZmVVVVZmZmVVVVZmZmVVVVVVVVZmZmVVVVZmZmZmZmZmZmd3d3d3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREVVVVREREVVVVVVVVZmZmVVVVZmZmVVVVZmZmVVVVZmZmd3d3d3d3d3d3iIiId3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmd3d3d3d3iIiId3d3ZmZmZmZmREREREREMzMzMzMzREREREREVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmVVVVVVVVZmZmd3d3d3d3d3d3ZmZmVVVVVVVVVVVVZmZmd3d3d3d3ZmZmVVVVVVVVVVVVREREVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVZmZmVVVVZmZmZmZmd3d3ZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREREREREREVVVVVVVVZmZmd3d3iIiIiIiImZmZmZmZiIiImZmZmZmZmZmZmZmZqqqqmZmZqqqqqqqqqqqqmZmZmZmZmZmZqqqqmZmZmZmZmZmZmZmZqqqqmZmZqqqqqqqqmZmZqqqqiIiImZmZiIiImZmZqqqqqqqqqqqqqqqqqqqqqqqqmZmZmZmZiIiIiIiImZmZmZmZmZmZmZmZmZmZqqqqmZmZqqqqqqqqqqqqqqqqqqqqqqqqu7u7qqqqqqqqqqqqqqqqqqqqqqqqqqqqu7u7u7u7zMzM7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u6qqqqqqqqqqqru7u6qqqru7u7u7u93d3d3d3bu7u8zMzMzMzN3d3d3d3e7u7t3d3d3d3czMzN3d3czMzN3d3czMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u6qqqru7u7u7u7u7u7u7u7u7u8zMzLu7u8zMzMzMzLu7u6qqqru7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqru7u6qqqru7u6qqqru7u7u7u6qqqpmZmZmZmZmZmYiIiIiIiHd3d4iIiJmZmaqqqru7u8zMzN3d3d3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////93d3bu7u6qqqt3d3d3d3bu7u6qqqszMzN3d3d3d3f///////////////////+7u7v///////////////////+7u7t3d3czMzLu7u7u7u6qqqru7u5mZmZmZmZmZmZmZmZmZmZmZmaqqqqqqqru7u7u7u5mZmZmZmZmZmbu7u6qqqru7u7u7u7u7u7u7u7u7u8zMzMzMzLu7u7u7u7u7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqru7u7u7u7u7u6qqqru7u6qqqru7u7u7u6qqqru7u6qqqru7u6qqqqqqqru7u7u7u8zMzLu7u6qqqoiIiGZmZlVVVURERERERDMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzMyIiIjMzMyIiIjMzMyIiIiIiIjMzMyIiIiIiIiIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIjMzMzMzM0RERERERERERERERERERFVVVVVVVVVVVVVVVURERERERERERERERERERERERERERDMzMzMzM0RERFVVVWZmZkRERDMzM0RERERERERERFVVVURERFVVVVVVVVVVVVVVVURERERERERERERERERERERERDMzM0RERERERERERERERFVVVURERFVVVVVVVVVVVWZmZlVVVVVVVVVVVURERERERERERERERDMzM1VVVVVVVVVVVVVVVWZmZnd3d2ZmZmZmZnd3d4iIiIiIiHd3d4iIiIiIiIiIiGZmZmZmZlVVVWZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZkRERDMzM0RERERERERERERERERERERERERERDMzM0RERERERERERGZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVTMzM0RERERERERERFVVVVVVVVVVVURERFVVVVVVVURERFVVVURERGZmZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVVVVVURERERERFVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d3d3d1VVVWZmZlVVVVVVVVVVVVVVVWZmZmZmZlVVVURERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZlVVVURERERERERERFVVVWZmZlVVVVVVVURERFVVVVVVVVVVVVVVVVVVVWZmZnd3d4iIiHd3d2ZmZlVVVURERERERERERERERERERERERERERERERFVVVWZmZlVVVVVVVWZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZlVVVURERERERERERERERERERERERERERERERERERERERERERERERGZmZmZmZlVVVURERERERERERDMzM0RERERERDMzMzMzM0RERFVVVVVVVURERERERERERERERERERDMzMyIiIjMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERERERERERERERDMzMzMzM0RERERERERERFVVVURERERERERERERERDMzM0RERDMzM0RERERERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERDMzM0RERFVVVVVVVURERERERERERERERERERERERERERFVVVWZmZnd3d2ZmZlVVVVVVVURERERERERERFVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERFVVVVVVVURERERERERERGZmZnd3d3d3d1VVVVVVVURERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERDMzM0RERFVVVWZmZmZmZnd3d2ZmZmZmZlVVVURERERERERERERERERERERERERERFVVVURERERERERERERERDMzM0RERERERERERERERERERFVVVWZmZlVVVVVVVVVVVVVVVWZmZlVVVVVVVWZmZlVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVURERFVVVURERFVVVURERFVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d3d3d2ZmZnd3d2ZmZmZmZmZmZmZmZnd3d2ZmZmZmZlVVVVVVVURERERERERERDMzMzMzM0RERERERFVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVURERERERFVVVWZmZnd3d3d3d2ZmZnd3d2ZmZmZmZmZmZlVVVYiIiJmZmXd3d2ZmZlVVVVVVVWZmZlVVVVVVVWZmZnd3d2ZmZlVVVVVVVURERFVVVURERFVVVWZmZlVVVWZmZmZmZmZmZnd3d2ZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZnd3d1VVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVXd3d3d3d4iIiIiIiJmZmZmZmaqqqqqqqqqqqpmZmaqqqqqqqqqqqpmZmaqqqpmZmaqqqpmZmYiIiJmZmZmZmZmZmZmZmaqqqqqqqqqqqqqqqqqqqpmZmZmZmaqqqru7u7u7u7u7u8zMzLu7u8zMzLu7u7u7u7u7u7u7u7u7u6qqqru7u8zMzMzMzMzMzLu7u7u7u8zMzLu7u7u7u6qqqqqqqqqqqpmZmZmZmZmZmZmZmaqqqpmZmaqqqru7u7u7u93d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7u7u7d3d3MzMzd3d3d3d3d3d3MzMzMzMy7u7u7u7vMzMy7u7u7u7u7u7u7u7vMzMzMzMzMzMzMzMzMzMzd3d3u7u7u7u7d3d3MzMzd3d3d3d3u7u7u7u7d3d3d3d3MzMzMzMzMzMzMzMzMzMzMzMy7u7vMzMy7u7uqqqqZmZmqqqq7u7u7u7u7u7u7u7u7u7vMzMzMzMzMzMy7u7u7u7u7u7u7u7uqqqqqqqqqqqqqqqqqqqqqqqq7u7u7u7u7u7uqqqq7u7u7u7vMzMy7u7u7u7uqqqqqqqqZmZmZmZmZmZmZmZmZmZmqqqqqqqq7u7vMzMzd3d3u7u7u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////u7u7MzMy7u7vd3d3d3d27u7uqqqq7u7u7u7vd3d3u7u7////////////////////////////////u7u7u7u7u7u7u7u7MzMy7u7vd3d3d3d3d3d3MzMzMzMzMzMy7u7vMzMy7u7u7u7vMzMy7u7u7u7uqqqq7u7u7u7uqqqqqqqqZmZmZmZmZmZmqqqqZmZmZmZmqqqqZmZmZmZmZmZmqqqqqqqq7u7u7u7u7u7vMzMy7u7vMzMy7u7u7u7u7u7vMzMy7u7u7u7u7u7vMzMzd3d3d3d3MzMzd3d3MzMy7u7uqqqqIiIhmZmZEREQzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzNEREQzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNEREQzMzNERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVEREREREREREREREQzMzMzMzMzMzMzMzNERERERERERERERERERERERERVVVVVVVVVVVVEREQzMzMzMzMzMzNEREQzMzNEREQzMzNEREQzMzNEREREREQzMzNERERERERERERERERERERVVVVmZmZVVVVVVVVERERERERERERERERERERERERERERERERmZmZVVVVVVVVVVVVVVVVmZmZmZmZ3d3dmZmZmZmZmZmZ3d3d3d3eIiIh3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZ3d3dmZmZVVVVERERERERERERERERERERERERERERERERERERERERERERVVVVVVVV3d3dmZmZVVVVVVVVVVVVmZmZVVVUzMzNERERERERERERVVVVmZmZVVVVERERVVVVERERVVVVVVVVVVVVmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZVVVVVVVVVVVVVVVVERERERERVVVVVVVVVVVVERERERERVVVVmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZVVVVVVVVmZmZmZmZVVVVERERERERERERERERERERVVVVERERVVVVERERVVVVERERVVVVmZmZ3d3d3d3d3d3d3d3dmZmZ3d3dmZmZVVVVERERERERERERVVVVmZmZVVVVVVVVERERVVVVERERVVVVVVVVVVVVmZmZ3d3d3d3dmZmZVVVVEREREREREREQzMzNERERERERERERERERVVVVVVVVVVVVERERERERVVVVmZmZ3d3dmZmZVVVVVVVVVVVVEREREREREREREREQzMzNEREREREREREQzMzNEREQzMzMzMzMzMzNERERERERVVVVmZmZmZmZVVVVERERERERERERERERVVVVmZmZmZmZmZmZVVVVEREREREQzMzNEREREREQzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzNERERVVVVEREREREQzMzMzMzMzMzMzMzNERERERERERERERERERERVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNERERERERVVVVERERVVVVVVVVERERERERERERVVVVmZmZERERERERERERERERERERERERERERVVVVVVVVVVVVEREREREREREREREREREQzMzMzMzMzMzMzMzNERERERERVVVVEREREREREREQzMzMzMzNERERmZmZ3d3d3d3dmZmZVVVVVVVVVVVVERERERERVVVVVVVVVVVVmZmZVVVVVVVVEREREREREREQzMzMzMzNERERERERVVVVVVVVVVVVmZmZVVVVVVVVEREREREQzMzNERERVVVVVVVVERERVVVVERERVVVVERERERERERERERERVVVVERERVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVERERERERVVVVERERERERERERERERVVVVVVVVEREREREQzMzNERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3dmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERERERERERVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVmZmZmZmZVVVVERERVVVVERERVVVVVVVVVVVVmZmZmZmZ3d3dmZmZVVVVmZmZmZmZmZmZmZmZ3d3eIiIhmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVV3d3d3d3dVVVVERERVVVVERERVVVVVVVVVVVVmZmZmZmZmZmZmZmZ3d3d3d3d3d3dmZmZmZmZVVVVVVVVVVVVmZmZVVVVERERVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3dmZmZmZmZmZmZVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3eIiIiZmZmqqqqZmZmqqqqZmZmqqqqqqqqqqqqqqqqqqqqZmZmZmZmZmZmZmZmqqqqZmZmqqqqqqqqqqqqqqqq7u7u7u7uqqqq7u7uqqqq7u7u7u7vMzMzd3d3d3d27u7vd3d3d3d3d3d3d3d3MzMzd3d3d3d3u7u7d3d3u7u7d3d3d3d3MzMyqqqqqqqqZmZmZmZmIiIiIiIiIiIiIiIiZmZmZmZmqqqqqqqrMzMzd3d3///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u3d3d3d3d7u7u3d3d7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzM3d3d3d3d7u7u7u7u7u7u3d3d3d3dzMzMzMzMu7u7u7u7u7u7u7u7u7u7qqqqu7u7u7u7u7u7zMzMu7u7zMzMu7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqqqqqqqqqu7u7qqqqu7u7u7u7u7u7zMzMu7u7u7u7u7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqqqqqqqqqzMzMzMzM3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7uzMzMu7u7zMzMu7u7qqqqqqqqqqqqu7u73d3d7u7u7u7u////////////////////////////////////7u7u3d3dzMzM3d3d3d3d3d3d3d3d3d3dzMzM3d3d3d3dzMzMzMzMu7u7u7u7u7u7qqqqmZmZiIiIiIiId3d3d3d3mZmZmZmZmZmZqqqqqqqqu7u7u7u7u7u7qqqqu7u7u7u7u7u7u7u7zMzMu7u7zMzMzMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMqqqqmZmZd3d3VVVVREREMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREREREREREREREVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREREREMzMzREREREREREREREREMzMzREREREREVVVVREREREREREREREREVVVVREREMzMzREREMzMzREREMzMzREREREREMzMzREREMzMzREREMzMzREREREREREREREREMzMzREREREREREREMzMzMzMzREREREREREREREREREREMzMzREREREREREREVVVVVVVVVVVVVVVVZmZmZmZmVVVVZmZmZmZmZmZmd3d3d3d3ZmZmVVVVZmZmd3d3d3d3d3d3d3d3ZmZmZmZmd3d3ZmZmZmZmVVVVREREREREREREMzMzREREREREREREMzMzREREVVVVVVVVZmZmVVVVVVVVREREVVVVVVVVZmZmVVVVMzMzREREVVVVVVVVVVVVVVVVREREVVVVREREVVVVVVVVVVVVVVVVd3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVREREREREREREREREREREREREVVVVREREREREREREVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVREREREREREREREREREREREREREREVVVVREREVVVVVVVVREREVVVVVVVVZmZmZmZmd3d3iIiId3d3ZmZmREREREREREREREREVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREZmZmd3d3d3d3VVVVREREREREREREREREREREREREREREVVVVREREREREREREREREREREMzMzREREVVVVVVVVZmZmZmZmZmZmREREREREVVVVREREREREMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREZmZmZmZmZmZmZmZmVVVVVVVVREREZmZmZmZmVVVVVVVVREREREREMzMzMzMzMzMzMzMzMzMzREREREREVVVVVVVVREREVVVVREREVVVVVVVVREREREREMzMzMzMzMzMzMzMzMzMzREREREREVVVVREREREREREREVVVVVVVVVVVVZmZmVVVVZmZmVVVVVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREREREVVVVVVVVVVVVVVVVREREMzMzMzMzMzMzREREMzMzMzMzREREREREREREVVVVVVVVZmZmZmZmZmZmVVVVREREREREMzMzREREREREREREVVVVREREREREREREMzMzREREMzMzMzMzVVVVZmZmd3d3d3d3ZmZmZmZmVVVVVVVVVVVVREREREREVVVVZmZmZmZmREREREREMzMzMzMzMzMzREREREREVVVVVVVVREREMzMzREREREREREREREREREREREREVVVVREREREREVVVVREREREREVVVVREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREVVVVREREREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVREREVVVVVVVVREREREREVVVVREREVVVVVVVVVVVVZmZmZmZmd3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREVVVVREREVVVVVVVVREREVVVVREREVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3ZmZmVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREREREVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVREREREREREREVVVVZmZmd3d3d3d3ZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmd3d3ZmZmVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmd3d3d3d3d3d3d3d3ZmZmZmZmVVVVVVVVZmZmd3d3ZmZmVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmd3d3d3d3d3d3d3d3iIiIiIiIZmZmZmZmd3d3d3d3d3d3d3d3d3d3iIiIiIiImZmZmZmZqqqqmZmZqqqqqqqqmZmZqqqqqqqqmZmZqqqqmZmZqqqqu7u7u7u7qqqqu7u7zMzMu7u7u7u7u7u7u7u7qqqqu7u7qqqqu7u7zMzMzMzMu7u7zMzM3d3d3d3dzMzMu7u7zMzMzMzMzMzMu7u7zMzMu7u7u7u7qqqqqqqqmZmZmZmZiIiIiIiIiIiIiIiImZmZmZmZqqqqu7u7zMzM7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3czMzN3d3d3d3d3d3czMzN3d3d3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzLu7u8zMzMzMzMzMzMzMzMzMzLu7u8zMzLu7u7u7u6qqqqqqqpmZmaqqqpmZmaqqqru7u6qqqru7u7u7u7u7u8zMzMzMzLu7u7u7u6qqqqqqqqqqqqqqqqqqqqqqqru7u7u7u8zMzMzMzN3d3d3d3e7u7v///+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7szMzLu7u7u7u5mZmYiIiJmZmaqqqru7u93d3e7u7u7u7v///////////+7u7v///////////+7u7t3d3czMzN3d3d3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3czMzMzMzLu7u7u7u8zMzLu7u8zMzLu7u6qqqqqqqru7u8zMzMzMzMzMzMzMzLu7u7u7u7u7u6qqqru7u7u7u8zMzMzMzMzMzMzMzN3d3d3d3d3d3d3d3e7u7t3d3e7u7u7u7t3d3d3d3d3d3czMzKqqqpmZmXd3d1VVVTMzMzMzMzMzMyIiIiIiIjMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzM0RERERERFVVVVVVVVVVVWZmZmZmZlVVVVVVVWZmZmZmZlVVVVVVVURERERERDMzMzMzMyIiIjMzMzMzMzMzM0RERDMzM0RERERERERERERERERERERERFVVVURERFVVVURERERERERERDMzM0RERFVVVURERERERERERERERERERERERERERERERFVVVVVVVURERERERERERFVVVURERFVVVURERERERERERFVVVURERERERERERERERDMzM0RERDMzM0RERDMzMzMzM0RERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVXd3d4iIiJmZmZmZmYiIiGZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVURERERERERERERERERERERERERERFVVVVVVVVVVVURERERERERERFVVVVVVVVVVVVVVVTMzM0RERFVVVVVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVWZmZnd3d3d3d3d3d2ZmZnd3d2ZmZlVVVWZmZmZmZlVVVVVVVURERERERERERFVVVVVVVVVVVURERFVVVURERERERFVVVVVVVVVVVWZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVURERERERERERDMzM0RERDMzM0RERERERERERFVVVURERFVVVURERFVVVVVVVWZmZoiIiHd3d3d3d1VVVURERFVVVURERERERERERFVVVURERERERERERERERERERERERERERFVVVWZmZnd3d3d3d1VVVVVVVURERERERDMzM0RERERERERERERERERERFVVVURERERERERERERERERERFVVVVVVVWZmZmZmZlVVVVVVVURERERERERERDMzM0RERERERDMzMzMzMzMzM0RERDMzM0RERERERDMzMzMzM0RERFVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZkRERERERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVWZmZlVVVVVVVVVVVVVVVTMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERDMzMzMzMzMzM0RERFVVVURERFVVVWZmZlVVVVVVVTMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzMzMzM0RERERERERERERERFVVVVVVVURERDMzMzMzMzMzMzMzMzMzM0RERERERERERERERFVVVVVVVWZmZmZmZmZmZmZmZlVVVURERERERERERERERERERERERERERERERERERDMzM0RERERERERERERERGZmZnd3d4iIiGZmZmZmZlVVVVVVVVVVVURERFVVVXd3d2ZmZlVVVVVVVURERERERCIiIjMzM0RERERERERERERERERERERERERERERERERERFVVVVVVVVVVVVVVVURERERERERERERERERERERERERERDMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERDMzM0RERERERERERFVVVVVVVURERFVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERFVVVVVVVVVVVWZmZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZlVVVURERFVVVURERERERERERERERERERERERERERERERFVVVURERERERERERDMzM0RERDMzM0RERERERERERDMzM0RERGZmZnd3d3d3d1VVVVVVVVVVVURERERERERERERERERERERERERERFVVVWZmZmZmZmZmZlVVVWZmZlVVVURERERERERERERERERERFVVVVVVVVVVVURERERERFVVVWZmZnd3d2ZmZlVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVXd3d2ZmZkRERERERFVVVVVVVURERFVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVURERERERFVVVURERFVVVVVVVVVVVWZmZoiIiHd3d4iIiHd3d3d3d2ZmZlVVVVVVVWZmZnd3d3d3d2ZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d4iIiIiIiHd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZnd3d4iIiHd3d3d3d3d3d2ZmZnd3d3d3d3d3d4iIiIiIiIiIiIiIiJmZmYiIiJmZmaqqqpmZmZmZmYiIiJmZmZmZmaqqqpmZmZmZmaqqqqqqqru7u6qqqru7u7u7u7u7u7u7u6qqqpmZmaqqqqqqqru7u6qqqqqqqru7u8zMzLu7u6qqqru7u8zMzLu7u7u7u6qqqqqqqpmZmZmZmZmZmaqqqpmZmaqqqpmZmZmZmYiIiIiIiIiIiIiIiIiIiJmZmbu7u8zMzN3d3f///////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3MzMzMzMzMzMzd3d3MzMzd3d3MzMzMzMzMzMzMzMzMzMzMzMzd3d3d3d3u7u7d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMy7u7u7u7u7u7uqqqqZmZmZmZmZmZmZmZmZmZmqqqqZmZmqqqqqqqq7u7u7u7u7u7u7u7u7u7vMzMy7u7u7u7u7u7u7u7u7u7vMzMzMzMzd3d3d3d3d3d3u7u7u7u7////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////u7u7d3d3d3d2qqqp3d3d3d3eZmZmqqqq7u7u7u7vMzMzMzMzd3d3////////////u7u7u7u7d3d3MzMzMzMzMzMzMzMzd3d3d3d3d3d3d3d3u7u7d3d3d3d3d3d3d3d3MzMzMzMzd3d3d3d3d3d3d3d3d3d3MzMzd3d3MzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7vMzMzd3d3MzMzd3d3MzMzd3d3MzMzMzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7uqqqqZmZmZmZmIiIiIiIhmZmZVVVVEREQzMzNEREQzMzNERERERERERERERERVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVERERVVVVEREREREREREREREQzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiJERERVVVUzMzMzMzMzMzNEREREREQzMzNERERERERERERVVVVVVVVERERERERERERERERERERERERERERVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNEREQzMzNEREREREREREREREREREREREREREREREQzMzMzMzNEREREREREREQzMzNERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVmZmaIiIiIiIiZmZlmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZVVVVVVVVERERERERERERERERmZmZmZmZVVVVmZmZVVVVVVVVERERERERERERVVVVVVVVVVVUzMzNERERERERERERERERERERERERVVVVERERERERVVVVVVVVmZmZmZmZ3d3dmZmZ3d3dmZmZVVVVVVVVmZmZ3d3dVVVVVVVVERERERERERERERERERERVVVVERERVVVVERERERERVVVVERERVVVVVVVVVVVVERERVVVVmZmZmZmZmZmZmZmaIiIh3d3dVVVVEREQzMzNERERERERERERERERERERERERERERERERERERERERERERERERVVVVmZmZ3d3d3d3dmZmZVVVVEREQzMzNERERERERERERVVVVEREREREREREQzMzNERERERERERERERERmZmZ3d3dmZmZVVVVEREREREREREREREREREQzMzNERERERERERERERERERERVVVVVVVVVVVVERERVVVVVVVVmZmZmZmZVVVVEREREREREREREREQzMzMzMzMzMzMzMzNERERVVVVVVVVEREREREREREQzMzMzMzMzMzNERERERERERERERERVVVVmZmZmZmZVVVVEREQzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzNERERERERERERmZmZVVVVmZmZVVVVEREREREQzMzMzMzMzMzMzMzNEREREREREREREREQzMzMzMzMzMzMzMzMzMzNERERERERVVVVVVVVEREQzMzMzMzMzMzMzMzMiIiIiIiIiIiIzMzNEREREREREREQzMzMzMzMzMzNERERERERERERVVVVVVVUzMzMzMzMiIiIzMzMzMzMzMzMiIiJERERERERVVVVERERERERVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVEREREREQzMzMzMzMzMzMzMzNERERERERVVVV3d3d3d3d3d3d3d3dmZmZmZmZmZmZ3d3dmZmZmZmZVVVVVVVVVVVVVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERERERVVVVVVVVEREREREQzMzNEREREREREREREREQzMzNEREQzMzNEREQzMzMzMzNERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVEREREREQzMzNEREREREREREREREQzMzMzMzMzMzMzMzNERERVVVV3d3d3d3eIiIh3d3d3d3d3d3dmZmZmZmZVVVVEREREREREREREREQzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREREREREREREREREREQzMzMzMzMzMzMzMzNERERERERERERERERVVVVmZmZ3d3dmZmZVVVVERERERERERERERERERERERERERERVVVV3d3d3d3dmZmZVVVVVVVVERERVVVVERERERERERERVVVVVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVmZmZERERVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVERERERERERERERERERERVVVVVVVVVVVVVVVVmZmZmZmZVVVVERERERERERERVVVVVVVVVVVVmZmZ3d3d3d3d3d3d3d3d3d3eIiIhmZmZVVVVmZmaIiIiIiIh3d3dmZmZVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3eIiIiIiIiIiIiIiIh3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3eIiIh3d3eIiIiIiIiZmZmIiIiZmZmZmZmIiIiZmZmZmZmqqqqqqqqqqqqZmZmZmZmqqqq7u7uqqqqZmZmZmZmIiIiZmZmqqqqqqqqqqqqqqqq7u7uqqqqZmZmZmZmZmZmqqqqqqqqqqqqqqqqqqqqZmZmIiIiZmZmZmZmZmZmIiIiIiIiIiIiIiIiZmZmZmZmZmZmZmZmqqqq7u7vd3d3u7u7////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////7u7u7u7u7u7u3d3d7u7u3d3d7u7u3d3d7u7u3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMu7u7u7u7qqqqqqqqu7u7u7u7qqqqmZmZmZmZqqqqmZmZmZmZqqqqqqqqqqqqqqqqu7u7u7u7zMzMzMzMzMzMzMzMzMzMzMzMzMzM3d3d3d3d7u7u7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3dzMzMqqqqd3d3d3d3mZmZqqqqu7u7u7u7u7u7u7u73d3d7u7u3d3dzMzMzMzMu7u7qqqqqqqqu7u7zMzMzMzM3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzMzMzMqqqqu7u7u7u7zMzMu7u7zMzMu7u7zMzMu7u7zMzMzMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7qqqqqqqqqqqqu7u7qqqqqqqqqqqqmZmZmZmZmZmZd3d3d3d3d3d3ZmZmZmZmZmZmZmZmd3d3ZmZmd3d3d3d3ZmZmZmZmZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzIiIiMzMzMzMzREREREREMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREREREREREREREVVVVREREVVVVVVVVVVVVVVVVREREREREMzMzREREREREREREREREREREREREREREREREREREVVVVREREREREREREREREREREREREVVVVREREREREVVVVVVVVZmZmVVVVZmZmZmZmVVVVZmZmZmZmd3d3iIiId3d3ZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmREREREREREREREREREREREREVVVVREREREREREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmd3d3d3d3VVVVVVVVREREVVVVREREREREVVVVREREREREREREREREREREREREVVVVREREVVVVREREVVVVVVVVZmZmZmZmVVVVd3d3iIiId3d3REREREREREREMzMzREREREREREREREREREREVVVVVVVVREREREREMzMzREREREREVVVVd3d3d3d3ZmZmVVVVREREREREMzMzREREREREREREREREREREREREMzMzMzMzREREREREREREZmZmd3d3VVVVREREREREREREREREREREMzMzREREMzMzREREVVVVREREREREREREVVVVREREREREREREVVVVZmZmZmZmVVVVREREREREMzMzREREMzMzMzMzREREREREVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREVVVVVVVVZmZmREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREREREREREREREVVVVZmZmVVVVVVVVMzMzMzMzMzMzMzMzMzMzMzMzMzMzVVVVREREREREREREREREMzMzMzMzMzMzREREREREVVVVVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzREREMzMzMzMzMzMzMzMzREREREREREREVVVVMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzREREVVVVREREREREVVVVZmZmZmZmVVVVVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREVVVVZmZmd3d3d3d3ZmZmZmZmZmZmd3d3iIiIVVVVVVVVVVVVREREREREREREVVVVREREMzMzMzMzIiIiIiIiMzMzMzMzMzMzREREREREREREREREREREREREVVVVVVVVMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzREREREREVVVVREREREREREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREREREZmZmd3d3d3d3d3d3ZmZmVVVVVVVVVVVVVVVVVVVVREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREVVVVVVVVREREREREREREREREREREREREREREREREVVVVVVVVREREVVVVZmZmZmZmVVVVVVVVVVVVREREREREVVVVREREREREVVVVVVVVd3d3ZmZmVVVVVVVVREREREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREVVVVVVVVZmZmVVVVREREREREVVVVREREVVVVVVVVVVVVVVVVREREVVVVZmZmZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmd3d3iIiId3d3iIiId3d3d3d3VVVVZmZmd3d3d3d3iIiId3d3ZmZmVVVVZmZmVVVVZmZmZmZmZmZmZmZmd3d3iIiId3d3iIiId3d3ZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3iIiId3d3iIiImZmZmZmZmZmZmZmZqqqqmZmZiIiIiIiIiIiImZmZiIiIiIiId3d3d3d3mZmZmZmZiIiIiIiImZmZiIiImZmZiIiIiIiImZmZmZmZmZmZmZmZmZmZqqqqmZmZmZmZmZmZmZmZiIiIiIiIiIiIiIiIiIiImZmZqqqqu7u73d3d3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u////////////////7u7u////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7t3d3d3d3d3d3d3d3e7u7t3d3d3d3d3d3czMzMzMzMzMzLu7u8zMzMzMzMzMzN3d3czMzMzMzMzMzMzMzLu7u8zMzLu7u7u7u6qqqqqqqqqqqqqqqqqqqqqqqru7u7u7u7u7u7u7u7u7u8zMzLu7u7u7u7u7u8zMzLu7u8zMzMzMzMzMzN3d3d3d3d3d3e7u7u7u7u7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7szMzKqqqpmZmYiIiJmZmaqqqru7u7u7u5mZmZmZmZmZmaqqqru7u6qqqqqqqru7u6qqqpmZmaqqqru7u7u7u8zMzMzMzMzMzMzMzMzMzN3d3d3d3d3d3czMzN3d3d3d3czMzMzMzLu7u8zMzLu7u7u7u7u7u7u7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqru7u7u7u8zMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u6qqqqqqqru7u6qqqru7u6qqqpmZmZmZmZmZmYiIiIiIiIiIiHd3d4iIiHd3d2ZmZmZmZmZmZmZmZnd3d2ZmZmZmZnd3d3d3d1VVVWZmZmZmZlVVVVVVVWZmZlVVVVVVVVVVVURERERERDMzM0RERDMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzM0RERDMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzM0RERDMzM0RERDMzM0RERFVVVVVVVVVVVURERERERERERERERERERERERFVVVURERERERDMzM0RERERERDMzM0RERERERERERFVVVURERERERERERFVVVURERFVVVURERFVVVURERERERERERERERERERERERFVVVURERERERERERFVVVVVVVWZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d4iIiHd3d3d3d3d3d2ZmZlVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVVVVVURERERERERERERERFVVVVVVVURERFVVVVVVVVVVVVVVVVVVVWZmZnd3d3d3d3d3d1VVVVVVVVVVVURERFVVVURERERERERERFVVVURERFVVVURERERERERERERERFVVVVVVVVVVVVVVVWZmZlVVVVVVVXd3d4iIiGZmZlVVVURERERERERERERERFVVVURERERERERERERERFVVVURERERERDMzMzMzMzMzM1VVVWZmZnd3d2ZmZkRERERERDMzM0RERDMzM0RERERERERERERERERERDMzM0RERDMzM0RERERERFVVVWZmZlVVVVVVVURERERERERERERERERERDMzM0RERERERERERERERERERFVVVVVVVURERDMzM0RERERERFVVVVVVVVVVVURERERERERERDMzMzMzMzMzM0RERERERERERERERDMzMyIiIjMzMzMzMzMzMzMzM0RERERERDMzM0RERFVVVWZmZlVVVURERDMzM0RERERERDMzMzMzMyIiIjMzM0RERDMzM0RERERERDMzM0RERDMzM0RERDMzM0RERERERGZmZlVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzM1VVVURERERERERERDMzMzMzMzMzMzMzM0RERERERERERERERERERDMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzM0RERDMzM0RERDMzMzMzMzMzM0RERERERERERFVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERFVVVURERERERERERFVVVWZmZlVVVURERERERERERERERERERDMzM0RERDMzMzMzM0RERERERERERFVVVXd3d3d3d3d3d2ZmZmZmZnd3d2ZmZlVVVVVVVURERDMzM0RERERERDMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERERERDMzM0RERFVVVVVVVURERFVVVURERERERERERDMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERFVVVVVVVURERERERERERFVVVVVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERFVVVVVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVURERERERFVVVVVVVVVVVTMzM0RERDMzM0RERERERERERDMzM0RERDMzM0RERERERERERFVVVVVVVVVVVVVVVTMzM0RERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERFVVVWZmZlVVVVVVVVVVVURERFVVVURERERERFVVVVVVVURERFVVVWZmZmZmZmZmZmZmZlVVVVVVVWZmZlVVVVVVVURERERERFVVVURERERERFVVVVVVVWZmZlVVVURERERERERERERERERERERERFVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d3d3d3d3d3d3d3d3d2ZmZmZmZlVVVXd3d3d3d3d3d4iIiHd3d2ZmZmZmZlVVVVVVVWZmZmZmZmZmZnd3d2ZmZnd3d3d3d3d3d2ZmZlVVVVVVVWZmZnd3d2ZmZnd3d2ZmZmZmZnd3d2ZmZmZmZmZmZmZmZnd3d4iIiGZmZmZmZnd3d2ZmZmZmZmZmZnd3d3d3d4iIiIiIiIiIiIiIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiHd3d3d3d4iIiIiIiJmZmZmZmZmZmYiIiIiIiHd3d4iIiJmZmZmZmZmZmYiIiIiIiIiIiJmZmaqqqqqqqqqqqt3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3d3d3MzMy7u7u7u7u7u7u7u7vMzMzMzMzMzMy7u7vMzMy7u7vMzMy7u7u7u7u7u7vMzMy7u7u7u7vMzMy7u7vMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7d3d3MzMy7u7uZmZmIiIiZmZmqqqqqqqp3d3dERERVVVVmZmaZmZmqqqqqqqqqqqqqqqqqqqqqqqqqqqq7u7u7u7u7u7vMzMzMzMzMzMzMzMzMzMzMzMzd3d3MzMy7u7u7u7u7u7uqqqqqqqq7u7u7u7u7u7uqqqqqqqqqqqqqqqqZmZmqqqqqqqqqqqq7u7u7u7u7u7u7u7u7u7u7u7u7u7uqqqq7u7u7u7u7u7uqqqqZmZmqqqqqqqqIiIiIiIiIiIh3d3dmZmZmZmZ3d3dmZmZmZmZVVVVmZmZ3d3d3d3dmZmZ3d3d3d3dmZmZ3d3dmZmZERERVVVVVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIzMzMiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERERERVVVVEREREREREREREREQzMzNEREREREREREQzMzMzMzNEREQzMzMzMzNEREREREREREREREREREQzMzNEREREREREREQzMzNEREQzMzNEREREREQzMzMzMzMzMzMzMzMzMzNERERERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZ3d3d3d3eIiIiZmZmIiIiIiIiIiIhmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERERERVVVV3d3d3d3dmZmZmZmZVVVVERERERERVVVVERERERERERERVVVVERERERERERERERERVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZ3d3dmZmZVVVVERERVVVVERERVVVVERERVVVVERERVVVVERERVVVVVVVVEREQzMzNEREQzMzNERER3d3d3d3dmZmZEREREREREREQzMzNEREQzMzNEREQzMzNEREREREREREQzMzNERERERERERERVVVVmZmZVVVVEREREREREREQzMzNEREQzMzNEREREREQzMzNERERERERERERERERVVVVVVVUzMzNERERERERVVVVmZmZEREREREQzMzMzMzMzMzMzMzNEREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNERERERERVVVVVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNEREQzMzMzMzNEREQzMzMzMzNERERERERVVVVEREQzMzMzMzMzMzNEREQiIiIzMzMzMzNEREQzMzNEREREREQzMzMzMzMzMzMzMzNEREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzNEREQzMzMzMzMzMzNEREQzMzNERERVVVVEREQzMzMiIiIiIiIzMzMiIiIzMzMiIiIzMzMzMzMzMzNERERERERERERERERERERERERERERVVVVVVVVVVVVVVVVEREREREREREQzMzNEREQzMzNEREQzMzNERERERERERERVVVVVVVVmZmZmZmZ3d3d3d3dmZmZmZmZmZmZVVVVEREREREQzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNERERERERERERERERVVVVVVVVVVVVEREREREQzMzMzMzMiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNVVVVmZmZ3d3d3d3dVVVVERERERERERERVVVUzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERVVVVERERERERERERERERERERVVVVERERVVVVEREREREQzMzNERERVVVVVVVVVVVVEREREREREREREREREREREREREREREREQzMzNERERVVVVVVVVmZmZVVVVVVVVVVVVERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVERERERERERERERERERERERERERERERERVVVVERERVVVVmZmZmZmZVVVVERERVVVVERERERERVVVVVVVVERERVVVVVVVVmZmZmZmZmZmZmZmZERERVVVVERERERERERERVVVVERERERERVVVVERERERERmZmZmZmZVVVVVVVVERERERERVVVVERERVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZVVVVVVVVmZmZmZmZ3d3d3d3eIiIh3d3d3d3dmZmZmZmZVVVV3d3eIiIh3d3d3d3eIiIh3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3dVVVVmZmZVVVVVVVVmZmZmZmZmZmZmZmZ3d3d3d3dmZmZmZmZmZmZ3d3d3d3dmZgD//wAAZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZoiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiHd3d3d3d3d3d4iIiIiIiIiIiHd3d4iIiHd3d3d3d4iIiIiIiIiIiIiIiJmZmaqqqru7u8zMzN3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7d3d3d3d3MzMzd3d3d3d3d3d3d3d3d3d3u7u7d3d3u7u7d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7////u7u7u7u7u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////d3d3MzMzMzMyqqqqZmZmZmZmZmZl3d3dVVVUzMzNERERVVVWIiIiIiIiZmZmqqqq7u7u7u7u7u7uqqqqqqqq7u7u7u7u7u7u7u7vMzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7vMzMy7u7uqqqqqqqqqqqqqqqqqqqqqqqqqqqq7u7uqqqqZmZmqqqqqqqqZmZmqqqqqqqqZmZmIiIiZmZmIiIh3d3eIiIh3d3d3d3dmZmZmZmZ3d3dmZmZ3d3d3d3d3d3dmZmZVVVVVVVVEREREREREREQzMzMzMzMzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIzMzMzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMzMzNEREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMiIiIzMzNERERERERERERERERVVVVmZmZVVVVVVVVEREREREREREREREQzMzMzMzNEREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzNEREQzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzNEREQzMzMzMzNERERVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmaIiIiIiIiIiIiIiIiIiIh3d3dmZmZmZmZmZmZmZmZVVVVmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVEREQzMzMzMzMzMzNERERERERERERVVVVVVVVVVVVVVVVVVVVERERERERVVVVERERERERERERERERERERERERERERERERERERERERVVVVERERERERVVVVERERERERVVVVERERVVVVVVVV3d3d3d3dVVVVERERERERERERERERVVVVERERERERERERVVVVERERERERERERERERVVVVERERERERmZmZ3d3dmZmZVVVUzMzMzMzMzMzMzMzNEREQzMzNEREREREREREREREREREQzMzMzMzMzMzNERERmZmZVVVVEREREREREREREREREREQzMzMzMzNEREREREQzMzNEREQzMzNERERERERERERERERERERERERVVVVmZmZVVVVEREQzMzNEREQzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzNEREREREREREQzMzNEREREREREREQzMzNERERERERVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNEREQzMzNEREQzMzMzMzMiIiIzMzMzMzNEREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNEREQzMzMzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVUzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNEREQzMzNERERVVVVVVVVVVVVVVVVEREREREQzMzMzMzMzMzMzMzMzMzNEREQzMzNERERERERERERVVVVmZmZmZmZmZmZ3d3dmZmZ3d3d3d3dVVVVEREQzMzNEREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREREREREREREREREREREREREREQzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNERERERER3d3dmZmZmZmZERERERERERERVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzNERERVVVVVVVVEREREREQzMzMzMzMiIiIzMzNERERERERERERVVVVEREQzMzMzMzMzMzMzMzNERERERERERERVVVVERERERERERERERERERERERERERERERERVVVVVVVVERERVVVVERERVVVVVVVVmZmZERERERERERERVVVVERERERERERERERERERERVVVVVVVVVVVVVVVUzMzNEREREREREREREREQzMzNVVVV3d3dVVVVVVVVmZmZmZmZVVVVVVVVERERERERERERERERVVVVVVVVVVVVmZmZVVVVmZmZmZmZVVVVVVVVVVVVERERERERVVVVERERERERERERERERVVVVVVVVVVVVmZmZmZmZmZmZVVVVERERVVVVERERVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZ3d3d3d3d3d3dmZmZmZmZmZmZVVVVVVVVmZmZ3d3eIiIiIiIiIiIh3d3d3d3dmZmZVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZ3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZ3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIh3d3d3d3dmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3eIiIiZmZmIiIiZmZmIiIiqqqqZmZm7u7vMzMzd3d3///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u7u7u////7u7u////////////////7u7u////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3dzMzMzMzMu7u7iIiIiIiImZmZiIiId3d3VVVVVVVVd3d3mZmZmZmZiIiImZmZu7u7qqqqqqqqqqqqu7u7zMzMzMzMu7u7u7u7u7u7zMzMu7u7zMzMu7u7zMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7qqqqqqqqqqqqqqqqmZmZqqqqmZmZiIiIiIiImZmZmZmZiIiImZmZiIiIiIiIiIiIiIiIiIiIiIiId3d3iIiImZmZiIiIiIiIiIiId3d3ZmZmZmZmVVVVMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzREREMzMzMzMzREREREREREREREREREREREREMzMzIiIiMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzREREREREREREREREREREVVVVREREVVVVREREREREREREREREREREREREREREREREMzMzREREMzMzREREMzMzMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREVVVVVVVVVVVVREREVVVVREREREREREREREREREREREREVVVVZmZmZmZmd3d3ZmZmd3d3d3d3ZmZmZmZmZmZmd3d3ZmZmZmZmZmZmVVVVVVVVVVVVREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREMzMzMzMzREREVVVVVVVVREREREREVVVVVVVVREREVVVVREREREREVVVVVVVVREREVVVVREREREREREREREREREREREREVVVVVVVVREREREREREREREREREREVVVVZmZmiIiIZmZmVVVVREREREREVVVVVVVVVVVVREREREREREREREREVVVVREREREREREREREREREREMzMzVVVVd3d3ZmZmREREMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREREREREREMzMzMzMzMzMzREREZmZmVVVVREREMzMzREREREREREREMzMzREREMzMzREREREREMzMzREREREREMzMzREREREREREREVVVVVVVVZmZmZmZmVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzMzMzMzMzREREREREMzMzMzMzMzMzREREREREVVVVVVVVMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREVVVVVVVVVVVVREREREREREREMzMzREREREREMzMzREREREREMzMzREREVVVVVVVVVVVVVVVVZmZmd3d3d3d3d3d3d3d3d3d3ZmZmREREREREREREREREREREREREMzMzREREMzMzREREMzMzREREMzMzREREREREREREREREREREVVVVVVVVREREREREIiIiIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzREREREREREREMzMzREREREREVVVVd3d3VVVVMzMzREREVVVVREREREREZmZmREREREREVVVVVVVVVVVVVVVVREREREREREREMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREVVVVREREREREMzMzMzMzMzMzMzMzREREMzMzVVVVREREVVVVREREREREVVVVREREREREVVVVVVVVREREREREREREREREREREREREZmZmVVVVREREREREREREVVVVREREREREREREREREREREVVVVVVVVZmZmVVVVREREMzMzREREMzMzMzMzREREVVVVZmZmVVVVREREZmZmZmZmZmZmVVVVREREVVVVREREREREREREZmZmVVVVVVVVZmZmVVVVZmZmZmZmVVVVREREVVVVVVVVREREREREVVVVREREREREREREVVVVZmZmZmZmZmZmZmZmREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVREREVVVVZmZmZmZmZmZmZmZmd3d3ZmZmd3d3d3d3d3d3d3d3ZmZmZmZmVVVVVVVVZmZmZmZmZmZmiIiImZmZiIiId3d3d3d3ZmZmZmZmVVVVZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmd3d3ZmZmZmZmVVVVREREVVVVVVVVVVVVZmZmZmZmd3d3d3d3d3d3d3d3ZmZmd3d3iIiImZmZiIiId3d3iIiId3d3ZmZmZmZmZmZmZmZmd3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiId3d3iIiIiIiIiIiImZmZiIiImZmZmZmZqqqqu7u7zMzM3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7t3d3czMzLu7u5mZmYiIiKqqqqqqqpmZmYiIiHd3d4iIiKqqqpmZmbu7u7u7u8zMzLu7u8zMzMzMzN3d3czMzMzMzN3d3czMzMzMzN3d3czMzN3d3d3d3d3d3d3d3czMzMzMzMzMzLu7u7u7u8zMzLu7u6qqqqqqqqqqqpmZmZmZmYiIiHd3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiJmZmYiIiIiIiIiIiJmZmYiIiJmZmZmZmYiIiJmZmZmZmYiIiHd3d2ZmZlVVVURERERERDMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMyIiIjMzMyIiIiIiIjMzMyIiIjMzMzMzM0RERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzM0RERDMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzM0RERERERFVVVVVVVURERDMzM0RERDMzM0RERDMzM0RERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERDMzM0RERDMzM0RERERERFVVVWZmZlVVVVVVVVVVVURERERERERERERERERERERERERERERERERERERERFVVVVVVVWZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVURERERERERERERERERERFVVVURERFVVVURERERERFVVVVVVVVVVVURERFVVVURERERERFVVVVVVVURERERERERERERERERERFVVVVVVVURERERERFVVVURERERERFVVVVVVVVVVVWZmZoiIiHd3d1VVVURERERERERERFVVVVVVVURERERERERERERERERERERERERERERERERERERERDMzM0RERHd3d2ZmZkRERERERDMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERERERDMzMzMzMzMzMzMzM1VVVWZmZkRERERERDMzM0RERDMzM0RERERERERERERERDMzM0RERERERERERDMzM0RERERERERERERERFVVVWZmZmZmZmZmZlVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERDMzM0RERERERDMzMzMzMzMzM1VVVURERFVVVURERDMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzM0RERDMzM0RERDMzMzMzMzMzMzMzM0RERERERERERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzM0RERDMzMzMzM0RERFVVVURERDMzMzMzMyIiIjMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERCIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVVVVVVVVVVVVVURERERERERERDMzM0RERERERDMzMzMzM0RERERERFVVVWZmZlVVVVVVVWZmZoiIiIiIiIiIiHd3d3d3d1VVVVVVVURERDMzM0RERERERERERERERERERDMzMzMzMzMzM0RERERERERERERERERERERERERERDMzM0RERFVVVURERERERCIiIjMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM1VVVWZmZnd3d1VVVURERERERFVVVVVVVURERFVVVVVVVURERFVVVWZmZmZmZkRERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVTMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERERERERERERERFVVVVVVVVVVVVVVVURERFVVVURERERERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVURERERERERERFVVVVVVVURERFVVVWZmZmZmZlVVVURERERERDMzM0RERERERFVVVVVVVVVVVVVVVURERGZmZnd3d2ZmZmZmZkRERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVURERERERERERERERERERFVVVURERFVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVURERFVVVVVVVVVVVVVVVXd3d3d3d2ZmZnd3d2ZmZnd3d2ZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZnd3d3d3d4iIiHd3d3d3d2ZmZmZmZmZmZmZmZlVVVWZmZmZmZnd3d3d3d3d3d2ZmZmZmZnd3d2ZmZlVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d3d3d2ZmZnd3d3d3d4iIiHd3d4iIiIiIiHd3d2ZmZmZmZlVVVVVVVWZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d4iIiIiIiIiIiIiIiIiIiJmZmZmZmZmZmZmZmZmZmbu7u93d3d3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////d3d3MzMy7u7uIiIiIiIiqqqrMzMy7u7uqqqqZmZmZmZmqqqq7u7vMzMzMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzMzMzMzMzMzMzMzMzMzMy7u7u7u7uqqqqqqqqZmZmZmZmIiIiIiIiIiIh3d3d3d3eIiIiIiIiIiIiZmZmZmZmIiIiIiIiZmZmIiIiIiIh3d3eIiIh3d3d3d3dmZmZmZmZmZmZVVVVVVVVEREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzNEREREREREREREREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzNERERERERERERERERVVVVmZmZVVVVVVVUzMzNEREREREREREREREREREREREQzMzNERERERERERERERERVVVVmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmaIiIiIiIiIiIiZmZmZmZlmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVEREREREQzMzNVVVVVVVVVVVVVVVVERERERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERERERVVVVVVVVVVVVERERERERERERERERVVVVmZmZmZmZmZmZmZmZ3d3d3d3dVVVVEREREREREREREREREREREREREREQzMzNEREREREREREREREREREQzMzNEREQzMzNERER3d3dmZmZVVVVEREQzMzMzMzMzMzMzMzMzMzNEREQzMzNEREREREQzMzMzMzMzMzMzMzMzMzNVVVVVVVVVVVVEREREREREREREREREREREREQzMzNEREQzMzMzMzMzMzMzMzNEREREREQzMzNERERERERVVVVVVVV3d3dVVVVERERVVVVEREQzMzMzMzMzMzMzMzNEREQzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzNEREREREQzMzMzMzNERERVVVVVVVVEREQzMzNEREQzMzNEREQzMzMzMzMzMzNEREREREQzMzMzMzNEREQzMzNEREQzMzMzMzMzMzNEREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzNERERVVVVVVVVVVVVEREQzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMiIiJEREQzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzNERERERERVVVVmZmZVVVVVVVUzMzNEREQzMzNEREQzMzMzMzNEREREREQzMzNERERERERVVVVVVVVVVVVVVVVmZmZ3d3eZmZmIiIh3d3d3d3dVVVVEREREREREREREREREREREREREREREREQzMzMzMzMzMzMzMzNEREREREREREQzMzNERERERERERERVVVVVVVVEREQzMzMzMzMzMzMiIiIzMzMiIiIzMzNEREQzMzNEREQzMzNEREQzMzNERERmZmaIiIhVVVVERERERERERERVVVVERERERERERERERERVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERVVVVVVVVEREQzMzMzMzMiIiIzMzMzMzMzMzNEREQzMzNERERERERVVVVVVVVVVVVVVVVVVVVERERVVVVEREQzMzMzMzNERERERERVVVVERERERERmZmZmZmZERERERERERERERERVVVVERERERERVVVVVVVVVVVVmZmZmZmZVVVVEREREREQzMzNVVVVVVVVERERVVVVVVVVmZmZVVVV3d3dmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVERERVVVVmZmZ3d3dmZmZVVVVmZmZVVVVVVVVVVVVERERVVVVVVVVERERERERVVVVmZmZmZmZmZmZmZmZERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZERERERERERERERERVVVVmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZVVVVVVVVmZmZ3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZVVVVVVVVmZmZVVVVmZmZ3d3d3d3dmZmZmZmZmZmZ3d3dmZmZVVVVVVVVERERmZmZmZmZ3d3d3d3d3d3dmZmZVVVVVVVV3d3d3d3dmZmaIiIiIiIh3d3dmZmZmZmZmZmZmZmZmZmZVVVVmZmZ3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZ3d3d3d3d3d3eIiIiZmZmZmZmIiIiIiIiIiIiZmZmqqqqZmZmZmZmqqqrMzMzd3d3///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////7u7uzMzMqqqqiIiImZmZqqqqzMzMzMzMu7u7qqqqqqqqqqqqu7u7zMzMzMzM3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzMzMzM3d3dzMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7qqqqqqqqmZmZu7u7u7u7qqqqmZmZqqqqiIiImZmZmZmZmZmZiIiIiIiId3d3ZmZmZmZmVVVVVVVVREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzREREREREREREREREVVVVREREREREREREVVVVREREREREREREREREVVVVVVVVVVVVVVVVREREVVVVREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzMzMzREREMzMzREREMzMzMzMzMzMzMzMzREREREREMzMzMzMzMzMzREREREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmVVVVd3d3d3d3d3d3d3d3mZmZiIiId3d3ZmZmZmZmZmZmZmZmd3d3ZmZmZmZmREREREREVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVVVVVVVVVVVVVREREREREMzMzREREZmZmd3d3ZmZmZmZmVVVVZmZmZmZmZmZmVVVVVVVVREREREREREREREREREREREREREREVVVVREREREREREREREREREREMzMzREREd3d3ZmZmZmZmREREMzMzREREMzMzMzMzMzMzMzMzREREMzMzREREREREMzMzMzMzMzMzMzMzREREZmZmVVVVREREREREREREREREREREREREMzMzREREREREMzMzREREREREREREMzMzREREREREREREREREZmZmVVVVVVVVREREREREMzMzMzMzREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREMzMzREREREREREREVVVVREREREREREREREREMzMzREREMzMzMzMzMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREREREVVVVZmZmVVVVREREMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzREREMzMzMzMzMzMzREREVVVVVVVVVVVVMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzREREREREREREVVVVZmZmVVVVVVVVREREMzMzREREREREMzMzREREMzMzREREREREREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmiIiId3d3d3d3d3d3VVVVREREREREMzMzREREMzMzREREREREMzMzMzMzMzMzMzMzMzMzREREREREMzMzREREMzMzREREREREVVVVVVVVVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVVVVVVVVVVVVVREREREREREREREREREREVVVVREREVVVVVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVVVVVVVVVREREMzMzIiIiMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREREREVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREREREREREREREREREVVVVZmZmVVVVREREREREREREREREREREREREVVVVVVVVZmZmZmZmVVVVVVVVVVVVREREREREREREREREVVVVZmZmZmZmZmZmREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmd3d3d3d3ZmZmVVVVVVVVZmZmZmZmVVVVVVVVVVVVREREREREREREVVVVVVVVZmZmVVVVVVVVREREREREREREVVVVREREVVVVVVVVZmZmVVVVMzMzREREREREREREREREVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmVVVVZmZmZmZmVVVVZmZmVVVVZmZmZmZmVVVVZmZmd3d3ZmZmVVVVZmZmZmZmZmZmVVVVZmZmZmZmd3d3iIiId3d3d3d3ZmZmZmZmVVVVZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmd3d3ZmZmd3d3d3d3ZmZmd3d3ZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiImZmZiIiImZmZmZmZqqqqu7u7u7u77u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////+7u7u7u7ru7u5mZmZmZmYiIiKqqqszMzN3d3d3d3czMzLu7u8zMzMzMzN3d3czMzMzMzN3d3d3d3czMzN3d3czMzN3d3d3d3d3d3d3d3d3d3czMzN3d3czMzMzMzMzMzLu7u8zMzLu7u7u7u8zMzLu7u6qqqqqqqpmZmZmZmYiIiHd3d2ZmZmZmZkRERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERFVVVWZmZlVVVVVVVWZmZnd3d3d3d3d3d2ZmZkRERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d2ZmZmZmZlVVVVVVVURERERERERERDMzMzMzMzMzMyIiIiIiIjMzMzMzMzMzMyIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMyIiIiIiIiIiIjMzMyIiIjMzMzMzMyIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMyIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERDMzMzMzM0RERERERERERERERERERERERERERERERERERERERERERERERERERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d2ZmZmZmZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZkRERERERGZmZmZmZoiIiJmZmYiIiGZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVURERFVVVURERFVVVWZmZnd3d1VVVURERERERDMzM0RERERERGZmZoiIiHd3d1VVVURERERERFVVVWZmZmZmZlVVVURERERERERERERERERERERERERERERERFVVVURERERERDMzM0RERERERFVVVXd3d3d3d2ZmZkRERERERDMzMzMzM0RERDMzMzMzM0RERDMzM0RERDMzMzMzM0RERDMzM0RERFVVVWZmZmZmZkRERERERERERERERERERERERERERERERERERDMzMzMzMzMzM0RERERERERERERERFVVVWZmZlVVVVVVVVVVVURERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERDMzMzMzM0RERERERERERGZmZlVVVURERERERERERDMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzM0RERERERFVVVURERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVWZmZlVVVVVVVURERERERDMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzM0RERDMzM0RERFVVVVVVVVVVVVVVVVVVVTMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIkRERFVVVURERFVVVWZmZmZmZlVVVVVVVVVVVURERERERERERERERDMzM0RERERERFVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d4iIiHd3d3d3d2ZmZlVVVURERERERDMzM0RERDMzMzMzMzMzM0RERDMzMzMzMzMzM0RERERERDMzM0RERERERERERERERFVVVURERERERERERERERERERERERERERDMzMzMzM0RERDMzMzMzMzMzMzMzM0RERDMzMzMzM0RERFVVVVVVVURERERERERERERERDMzM0RERERERERERFVVVURERERERERERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVVVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERFVVVVVVVVVVVWZmZkRERFVVVURERERERERERERERERERERERFVVVWZmZlVVVVVVVWZmZmZmZlVVVVVVVURERFVVVURERGZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERFVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVURERERERERERFVVVXd3d1VVVVVVVURERERERERERERERFVVVVVVVVVVVWZmZmZmZlVVVURERERERERERFVVVURERFVVVVVVVWZmZmZmZmZmZnd3d3d3d3d3d3d3d2ZmZlVVVWZmZnd3d2ZmZmZmZmZmZnd3d3d3d3d3d1VVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVURERGZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVXd3d4iIiIiIiIiIiHd3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZnd3d2ZmZnd3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiJmZmZmZmZmZmaqqqru7u8zMzMzMzN3d3f///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////u7u67u7uqqqqIiIiIiIiqqqrd3d3////u7u7u7u7d3d3d3d3u7u7d3d3d3d3d3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3MzMzMzMy7u7u7u7uZmZmZmZmZmZmIiIhmZmZ3d3dmZmZVVVVVVVVVVVUzMzNEREQzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNVVVVERERVVVVERERVVVVVVVVmZmZmZmZmZmZmZmaIiIh3d3d3d3d3d3dmZmZ3d3d3d3dmZmZmZmZVVVVmZmZ3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZVVVVEREREREQzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIzMzMiIiIiIiIiIiIzMzMzMzMzMzMzMzMiIiIiIiIiIiIzMzMiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNEREQzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzNEREREREREREREREQzMzNEREQzMzNERERERERERERERERERERERERERERERERVVVVVVVVERERVVVVVVVVVVVVERERVVVVVVVVERERVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZVVVVERERERERmZmZ3d3d3d3eZmZmIiIh3d3d3d3dmZmZmZmZVVVVmZmZVVVVVVVVVVVVmZmZmZmZVVVVVVVVmZmZmZmZ3d3dmZmZVVVVVVVVERERVVVVVVVVmZmZ3d3d3d3dVVVVEREQzMzMzMzNVVVVmZmZmZmZmZmZVVVVEREQzMzNEREREREREREREREREREREREREREREREREREQzMzNERERmZmZ3d3dVVVVVVVVVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERERERERERVVVVmZmZmZmZERERERERERERERERERERERERVVVVERERERERERERERERERERERERERERVVVVmZmZmZmZVVVVERERERERVVVVmZmZVVVVEREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERmZmZVVVVVVVVEREREREQzMzNEREQzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVERERERERVVVVVVVVEREQzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVVVVVmZmZVVVVmZmZmZmZVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERmZmZmZmZVVVVVVVVVVVVVVVVEREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERERERERERVVVVVVVVVVVVmZmZ3d3d3d3eIiIiIiIiIiIh3d3dmZmZmZmZmZmZVVVVVVVVEREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzNERERERERVVVVERERERERERERERERVVVUzMzNERERERERVVVVEREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzNERERERERERERVVVVVVVVEREREREQzMzMzMzNEREQzMzMzMzNERERERERVVVVERERERERVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNERERVVVVVVVVmZmZmZmZVVVVEREREREQzMzNERERERERERERVVVVmZmZVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVmZmZVVVVmZmZVVVVmZmZVVVVVVVVEREREREQzMzNERERVVVVVVVVmZmZmZmZmZmZVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZVVVVVVVVVVVV3d3d3d3dVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVERERERERERERERERVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3dmZmZmZmZVVVVVVVVmZmZmZmZVVVVVVVVmZmZmZmZmZmZVVVVERERVVVVVVVVVVVVVVVVERERERERERERERERmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZ3d3eIiIh3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZmZmZmZmaIiIiIiIh3d3d3d3eIiIiIiIiIiIiZmZmZmZmZmZmqqqqZmZmqqqq7u7vMzMzMzMzu7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u////////////////////7u7u////////////////////////////////////7u7u3d3dqqqqiIiImZmZqqqq3d3d7u7u////7u7u7u7uzMzMu7u73d3d3d3d3d3d3d3d3d3d3d3d7u7uzMzMu7u7u7u7u7u7qqqqqqqqu7u7qqqqmZmZmZmZiIiIZmZmVVVVVVVVREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzREREREREMzMzREREMzMzMzMzREREVVVVVVVVVVVVZmZmZmZmd3d3d3d3ZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3iIiIiIiId3d3ZmZmd3d3d3d3d3d3d3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVREREMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzMzMzMzMzREREREREREREREREREREREREREREVVVVREREREREVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREVVVVVVVVVVVVVVVVREREVVVVREREVVVVVVVVREREVVVVZmZmd3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiId3d3ZmZmZmZmZmZmZmZmd3d3d3d3ZmZmVVVVZmZmd3d3d3d3ZmZmZmZmVVVVZmZmVVVVVVVVZmZmVVVVd3d3VVVVREREREREREREVVVVVVVVZmZmZmZmd3d3ZmZmVVVVREREREREREREREREREREREREREREREREREREREREREREVVVVd3d3ZmZmREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzREREVVVVZmZmd3d3ZmZmVVVVVVVVREREREREREREREREREREREREVVVVREREREREMzMzREREREREREREREREVVVVVVVVREREREREREREREREZmZmVVVVVVVVREREREREMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVZmZmZmZmZmZmVVVVZmZmVVVVREREREREREREMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVVVVVVVVVVVVVZmZmVVVVREREREREMzMzREREMzMzREREMzMzMzMzREREREREMzMzREREVVVVZmZmZmZmVVVVREREVVVVVVVVVVVVZmZmVVVVREREREREREREREREMzMzREREREREREREVVVVZmZmiIiIZmZmREREREREREREREREREREVVVVREREREREMzMzMzMzMzMzMzMzMzMzREREMzMzREREVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVZmZmVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVd3d3iIiImZmZmZmZiIiId3d3ZmZmZmZmZmZmREREVVVVREREVVVVVVVVREREREREREREMzMzMzMzMzMzMzMzMzMzREREREREVVVVVVVVVVVVREREREREMzMzMzMzMzMzREREVVVVVVVVVVVVREREMzMzREREMzMzREREMzMzREREMzMzREREVVVVVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVVVVVZmZmVVVVREREREREREREREREREREREREREREREREVVVVREREVVVVVVVVREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREVVVVVVVVZmZmZmZmVVVVVVVVREREREREVVVVREREVVVVVVVVZmZmZmZmVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmVVVVVVVVREREREREREREVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmVVVVVVVVREREMzMzREREREREREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVZmZmZmZmVVVVZmZmd3d3VVVVREREREREVVVVVVVVVVVVREREREREVVVVVVVVVVVVZmZmZmZmVVVVVVVVREREVVVVVVVVREREVVVVZmZmZmZmZmZmd3d3d3d3ZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVZmZmZmZmVVVVREREMzMzREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmd3d3d3d3iIiId3d3d3d3ZmZmZmZmd3d3ZmZmd3d3ZmZmZmZmVVVVd3d3ZmZmd3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiImZmZmZmZqqqqu7u7u7u7u7u7zMzM3d3d3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////93d3czMzO7u7u7u7v///////////////+7u7u7u7u7u7u7u7u7u7u7u7v///+7u7v///////////93d3bu7u5mZmYiIiIiIiKqqqru7u7u7u6qqqoiIiHd3d5mZmbu7u8zMzN3d3d3d3czMzMzMzKqqqqqqqru7u6qqqqqqqqqqqru7u6qqqqqqqpmZmYiIiHd3d1VVVURERERERERERDMzM0RERDMzM0RERDMzMzMzMzMzM0RERDMzM0RERERERERERFVVVVVVVVVVVWZmZmZmZlVVVWZmZmZmZlVVVWZmZoiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiHd3d4iIiIiIiHd3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVVVVVURERERERDMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIjMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIjMzMyIiIjMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERDMzM0RERDMzM0RERERERERERERERFVVVURERFVVVURERERERERERFVVVURERERERFVVVVVVVURERERERERERERERERERERERFVVVURERFVVVURERFVVVURERERERERERFVVVURERFVVVXd3d4iIiIiIiHd3d2ZmZnd3d3d3d3d3d4iIiHd3d3d3d2ZmZnd3d3d3d4iIiIiIiGZmZlVVVURERFVVVWZmZnd3d3d3d3d3d2ZmZlVVVVVVVURERFVVVVVVVWZmZlVVVURERFVVVVVVVVVVVVVVVVVVVVVVVXd3d2ZmZmZmZlVVVURERFVVVURERERERERERFVVVURERERERERERGZmZnd3d2ZmZkRERERERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERFVVVWZmZmZmZmZmZlVVVURERERERERERERERERERERERERERERERERERERERERERDMzMzMzM0RERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVURERFVVVURERERERERERDMzMzMzMzMzMzMzM0RERERERDMzM0RERERERFVVVWZmZnd3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVURERERERERERERERERERERERERERERERDMzM0RERDMzM0RERERERFVVVVVVVVVVVWZmZmZmZmZmZmZmZkRERERERERERERERERERERERDMzM0RERERERERERFVVVXd3d2ZmZlVVVVVVVURERERERFVVVVVVVVVVVWZmZlVVVVVVVURERERERERERERERERERFVVVXd3d2ZmZmZmZlVVVURERERERERERERERFVVVVVVVVVVVVVVVURERERERERERERERERERERERFVVVVVVVVVVVVVVVURERERERERERERERGZmZmZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVURERFVVVXd3d5mZmZmZmXd3d2ZmZmZmZlVVVURERFVVVURERERERFVVVVVVVVVVVURERERERERERERERERERERERERERERERDMzM1VVVVVVVVVVVURERERERDMzMzMzMzMzM0RERDMzM1VVVVVVVVVVVURERFVVVURERERERERERDMzM0RERERERFVVVVVVVVVVVURERDMzMzMzM0RERDMzM0RERDMzMzMzM0RERDMzM1VVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVURERFVVVURERERERERERERERERERFVVVURERERERERERDMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERFVVVVVVVVVVVWZmZnd3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZlVVVURERERERERERFVVVVVVVVVVVVVVVVVVVVVVVXd3d2ZmZlVVVURERERERERERERERERERFVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d1VVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d1VVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVWZmZlVVVURERFVVVVVVVVVVVWZmZlVVVVVVVWZmZnd3d2ZmZlVVVWZmZlVVVWZmZlVVVWZmZmZmZmZmZlVVVVVVVURERERERERERERERERERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVWZmZlVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZnd3d2ZmZmZmZnd3d2ZmZmZmZnd3d3d3d3d3d4iIiIiIiIiIiIiIiJmZmZmZmZmZmZmZmZmZmbu7u6qqqru7u7u7u8zMzMzMzO7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7MzMy7u7vMzMzu7u7d3d3d3d3MzMzd3d3MzMzMzMzMzMzd3d3u7u7u7u7u7u7u7u7////////////u7u7MzMyZmZlmZmZmZmZmZmZmZmZ3d3dmZmZmZmZ3d3eIiIiqqqq7u7uqqqqqqqqqqqqqqqqqqqq7u7vMzMy7u7vMzMy7u7u7u7u7u7uqqqqqqqqIiIh3d3dmZmZVVVVERERVVVVVVVVERERVVVVVVVVmZmZVVVVmZmZmZmZ3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIh3d3d3d3eIiIh3d3eIiIiZmZmIiIiIiIiIiIh3d3eIiIiIiIiIiIiIiIiIiIh3d3dmZmZmZmZmZmZVVVVVVVVVVVVEREQzMzNEREQzMzMzMzMzMzMiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIiIiIiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVEREREREREREQzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzNEREQzMzNEREQzMzMzMzMiIiIiIiIzMzMzMzMzMzMzMzNERERERERERERERERERERERERERERERERVVVVVVVVERERERERERERVVVVEREQzMzNEREREREREREQzMzNERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZmZmZ3d3d3d3dmZmZmZmZ3d3d3d3eIiIh3d3dVVVVERERERERERERERER3d3d3d3d3d3d3d3dVVVVmZmZERERERERVVVVmZmZ3d3dVVVVVVVVmZmZVVVVERERVVVVVVVVVVVVmZmZ3d3dmZmZmZmZVVVVERERERERERERERERERERERERERERERER3d3dmZmZVVVVEREREREREREREREREREREREREREREREQzMzMzMzMzMzNEREREREQzMzNVVVVmZmZmZmZmZmZVVVVVVVVVVVVERERERERVVVVEREREREQzMzNEREREREREREREREQzMzNERERERERERERERERERERERERERERmZmZVVVVERERERERERERVVVVERERVVVVVVVVVVVVEREQzMzNEREQzMzNEREQzMzMzMzNERERERERVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVERERVVVVVVVVVVVVERERVVVVERERERERERERERERERERERERERERERERERERERERERERVVVVmZmZ3d3dmZmZmZmZmZmZVVVVVVVVERERERERERERERERERERERERERERVVVV3d3d3d3dmZmZVVVVERERERERERERERERERERVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVmZmZmZmZ3d3dVVVVEREQzMzNEREQzMzMzMzNERERERERVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVERERERERERERERERERERVVVVmZmZVVVVmZmZmZmZVVVVmZmZVVVVVVVVVVVVmZmaIiIiIiIiIiIh3d3dmZmZVVVVmZmZVVVVERERERERERERERERVVVVVVVVmZmZVVVVERERERERERERERERERERERERERERVVVVVVVVVVVVEREREREREREQzMzNERERERERERERERERERERERERVVVVVVVVVVVVERERERERERERERERERERERERVVVVVVVVEREQzMzNEREQzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzNERERmZmZVVVVVVVVmZmZVVVVmZmZVVVVVVVVVVVVERERERERERERERERERERVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3dVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVERERVVVVERERVVVVVVVVmZmZVVVVERERERERERERERERERERERERVVVVVVVVmZmZmZmZVVVV3d3dmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3d3d3dmZmZ3d3dmZmZVVVVVVVVVVVVVVVVVVVVERERERERVVVVERERVVVVVVVVVVVVVVVVmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVmZmZVVVVmZmZmZmZmZmZVVVVERERERERERERERERERERVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZmZmZmZmZ3d3dmZmZmZmZ3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3d3d3dmZmZ3d3d3d3eIiIiIiIiIiIh3d3eIiIiIiIiZmZmZmZmZmZmqqqrMzMzMzMzMzMzd3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3diIiId3d3iIiIiIiId3d3iIiIiIiImZmZqqqqqqqqqqqqqqqqu7u7zMzMzMzM3d3dzMzM3d3d7u7u7u7uzMzMqqqqd3d3d3d3mZmZmZmZmZmZiIiId3d3d3d3d3d3iIiIiIiIiIiId3d3iIiImZmZmZmZmZmZqqqqqqqqqqqqu7u7qqqqqqqqqqqqqqqqmZmZmZmZiIiIiIiImZmZmZmZiIiIiIiImZmZiIiIiIiImZmZmZmZiIiIiIiImZmZiIiId3d3iIiIiIiIiIiId3d3mZmZmZmZiIiIiIiIiIiIiIiImZmZiIiId3d3iIiIiIiIZmZmVVVVZmZmVVVVREREREREREREMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVZmZmVVVVREREREREREREREREREREMzMzREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREMzMzMzMzMzMzREREMzMzREREREREREREMzMzREREREREVVVVMzMzMzMzMzMzMzMzREREMzMzREREREREREREVVVVVVVVVVVVVVVVVVVVREREREREVVVVREREREREMzMzREREVVVVREREREREVVVVd3d3ZmZmZmZmVVVVVVVVZmZmd3d3ZmZmZmZmZmZmVVVVREREREREMzMzMzMzREREd3d3iIiId3d3d3d3ZmZmVVVVVVVVREREVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVd3d3d3d3ZmZmZmZmd3d3ZmZmZmZmVVVVREREREREREREVVVVREREREREVVVVZmZmVVVVREREMzMzMzMzREREVVVVREREREREREREVVVVREREREREREREREREREREREREZmZmd3d3ZmZmREREMzMzVVVVVVVVVVVVVVVVREREREREREREREREREREREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVREREREREMzMzMzMzREREREREVVVVVVVVVVVVVVVVREREVVVVREREREREREREREREVVVVVVVVZmZmZmZmZmZmREREVVVVREREREREREREREREVVVVVVVVVVVVREREVVVVVVVVREREREREREREREREREREREREREREMzMzVVVVZmZmd3d3d3d3VVVVVVVVVVVVREREVVVVZmZmVVVVZmZmVVVVVVVVVVVVREREZmZmZmZmVVVVREREVVVVREREREREREREREREREREREREREREVVVVZmZmd3d3d3d3d3d3d3d3ZmZmZmZmREREREREMzMzMzMzMzMzREREMzMzMzMzMzMzREREREREVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREREREREREMzMzMzMzMzMzREREVVVVREREVVVVVVVVZmZmZmZmd3d3ZmZmZmZmd3d3d3d3d3d3d3d3VVVVVVVVREREREREREREREREREREREREREREREREVVVVVVVVZmZmZmZmVVVVREREREREVVVVREREREREVVVVVVVVREREREREREREMzMzREREMzMzREREREREREREMzMzREREVVVVZmZmVVVVVVVVREREREREREREREREVVVVREREREREMzMzMzMzREREMzMzREREMzMzMzMzMzMzMzMzMzMzREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVREREREREMzMzREREREREREREREREREREVVVVREREREREREREREREREREREREREREREREVVVVVVVVVVVVZmZmREREVVVVZmZmd3d3d3d3d3d3d3d3ZmZmVVVVVVVVREREREREVVVVVVVVZmZmZmZmZmZmVVVVVVVVREREVVVVREREVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREVVVVVVVVZmZmVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVZmZmZmZmZmZmd3d3ZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3d3d3d3d3ZmZmZmZmd3d3ZmZmVVVVVVVVVVVVREREVVVVVVVVREREREREVVVVZmZmZmZmVVVVVVVVZmZmVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmVVVVREREVVVVZmZmZmZmZmZmVVVVVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmd3d3d3d3d3d3d3d3d3d3ZmZmZmZmd3d3d3d3d3d3d3d3iIiIiIiImZmZiIiIiIiIiIiImZmZiIiImZmZqqqqu7u73d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7u7u7t3d3d3d3bu7u4iIiGZmZmZmZlVVVVVVVXd3d3d3d4iIiKqqqru7u6qqqqqqqpmZmbu7u8zMzLu7u5mZmZmZmbu7u8zMzN3d3czMzLu7u7u7u8zMzLu7u7u7u6qqqqqqqqqqqqqqqpmZmZmZmZmZmZmZmZmZmZmZmZmZmaqqqqqqqqqqqru7u7u7u7u7u7u7u7u7u8zMzMzMzLu7u6qqqqqqqqqqqpmZmZmZmYiIiJmZmZmZmXd3d4iIiJmZmYiIiIiIiIiIiHd3d3d3d4iIiJmZmZmZmZmZmZmZmZmZmYiIiIiIiIiIiIiIiHd3d2ZmZlVVVVVVVURERDMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERDMzMzMzMzMzM0RERERERERERERERDMzMyIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERERERERERDMzM0RERERERDMzM0RERDMzMzMzM0RERDMzMzMzMzMzMyIiIjMzMyIiIhERESIiIhERESIiIhERESIiIjMzMzMzMzMzMzMzM0RERDMzM0RERERERERERDMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERDMzMzMzM0RERERERERERERERFVVVVVVVURERFVVVURERFVVVURERERERERERFVVVURERFVVVURERDMzM1VVVWZmZlVVVURERFVVVVVVVVVVVURERERERFVVVURERFVVVURERFVVVURERERERDMzMzMzM0RERERERFVVVWZmZnd3d2ZmZnd3d1VVVVVVVWZmZkRERFVVVWZmZmZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZnd3d2ZmZlVVVVVVVURERFVVVURERGZmZmZmZmZmZkRERERERDMzM0RERERERERERERERERERERERERERFVVVURERDMzM0RERERERFVVVWZmZlVVVVVVVURERERERERERFVVVURERFVVVURERERERERERERERERERFVVVURERERERFVVVVVVVURERFVVVURERGZmZmZmZlVVVURERERERERERERERERERDMzM0RERDMzM0RERFVVVVVVVWZmZmZmZlVVVVVVVVVVVURERERERFVVVWZmZmZmZlVVVVVVVVVVVURERERERERERFVVVURERERERFVVVVVVVVVVVVVVVURERFVVVURERERERERERERERFVVVURERERERFVVVWZmZmZmZmZmZlVVVURERERERERERFVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZlVVVURERERERERERDMzM0RERDMzM0RERDMzMzMzM0RERGZmZmZmZmZmZmZmZnd3d2ZmZlVVVURERDMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERFVVVVVVVWZmZmZmZmZmZnd3d1VVVURERERERERERDMzM0RERDMzMzMzMzMzM1VVVURERFVVVVVVVWZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZlVVVURERERERERERERERERERERERERERERERDMzM0RERERERERERFVVVWZmZmZmZlVVVURERERERFVVVVVVVVVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERFVVVVVVVVVVVVVVVVVVVURERFVVVURERFVVVURERERERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERFVVVVVVVURERERERDMzM0RERERERDMzM0RERERERERERERERERERFVVVVVVVURERERERERERERERERERGZmZlVVVWZmZmZmZlVVVVVVVVVVVWZmZoiIiHd3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVURERFVVVVVVVURERFVVVVVVVWZmZmZmZlVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVURERFVVVXd3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d2ZmZnd3d3d3d3d3d1VVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d3d3d2ZmZmZmZmZmZmZmZmZmZnd3d2ZmZlVVVURERFVVVURERERERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVURERFVVVURERFVVVURERFVVVURERFVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d4iIiIiIiHd3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiJmZmYiIiJmZmZmZmbu7u7u7u8zMzN3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3MzMzMzMyqqqqZmZmZmZmIiIh3d3d3d3eIiIiZmZmqqqqqqqq7u7u7u7u7u7uqqqqqqqqZmZmIiIiZmZmqqqq7u7vMzMzMzMzMzMzMzMzMzMzMzMy7u7vMzMzMzMzMzMy7u7u7u7u7u7vMzMzMzMzMzMy7u7u7u7u7u7vMzMy7u7vMzMy7u7u7u7u7u7vMzMzMzMy7u7u7u7u7u7uZmZmqqqqZmZmIiIiZmZmIiIiZmZmZmZmIiIiZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmqqqqZmZmIiIh3d3d3d3dmZmZmZmZVVVVVVVVEREREREQzMzMzMzMzMzMzMzMiIiIiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMiIiIzMzMzMzNEREQzMzMzMzNEREREREQzMzNERERVVVVEREREREREREQzMzNEREQzMzNEREQzMzNEREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIiIiIzMzMiIiIiIiIiIiIREREiIiIREREiIiIREREREREREREiIiIzMzMiIiIzMzMzMzMzMzNEREREREQzMzNEREREREREREQzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNEREQzMzNEREQzMzNEREREREQzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzNERERERERERERERERVVVVVVVVERERERERERERVVVVERERVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVERERERERVVVVEREREREREREREREREREREREREREREREREREQzMzNEREQzMzMzMzNVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVERERVVVVmZmZVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZ3d3dmZmZmZmZVVVVVVVVVVVVmZmZmZmZmZmZEREREREREREREREQzMzNERERERERERERERERERERERERVVVVERERERERERERERERVVVVVVVVERERERERERERERERERERVVVVERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZVVVVERERERERERERERERERERERERERERERERERERVVVVVVVVVVVVmZmZ3d3dmZmZmZmZVVVVVVVVmZmZmZmZVVVVVVVVmZmZVVVVVVVVEREREREREREQzMzMzMzNERERVVVVVVVVVVVVERERVVVVERERERERERERERERERERERERERERVVVVmZmZmZmZmZmZVVVVERERERERERERERERVVVVERERVVVVVVVVmZmZmZmZmZmZ3d3dVVVVEREREREQzMzMzMzNEREQzMzNERERERERERERVVVVVVVVVVVVVVVVmZmZmZmZ3d3dmZmZEREQzMzNEREQzMzNEREQzMzMzMzMzMzNEREREREQzMzNERERVVVVVVVVVVVVmZmZ3d3dmZmZVVVUzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVEREREREREREREREQzMzMzMzMzMzNEREQzMzNERERERERERERERERVVVVmZmZVVVVVVVVVVVVVVVVmZmZVVVVEREREREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVEREQzMzNEREQzMzNEREQzMzMzMzMzMzMzMzMzMzNEREQzMzNERERERERVVVVERERVVVVVVVVEREREREQzMzNEREQzMzNEREREREQzMzNERERERERERERERERVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZ3d3d3d3d3d3dmZmZmZmZ3d3d3d3dmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZVVVVERERVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZVVVVVVVVVVVVERERVVVVVVVVVVVV3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZ3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZVVVVVVVVERERERERERERERERERERERERVVVVVVVVVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVERERERERERERVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVmZmZmZmZ3d3dmZmZVVVVVVVVmZmZmZmZ3d3d3d3eZmZmIiIiIiIh3d3eIiIiZmZmIiIiZmZmZmZmIiIiZmZmZmZm7u7vMzMzd3d3u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u////7u7u7u7uu7u7mZmZqqqqzMzMu7u7qqqqmZmZu7u7u7u7mZmZiIiIiIiIiIiIiIiImZmZqqqqqqqqqqqqqqqqqqqqu7u7qqqqqqqqqqqqqqqqmZmZmZmZmZmZqqqqqqqqqqqqu7u7zMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7zMzMu7u7u7u7u7u7u7u7qqqqqqqqu7u7u7u7mZmZqqqqu7u7qqqqqqqqqqqqmZmZmZmZiIiIiIiIiIiIZmZmZmZmZmZmVVVVREREREREMzMzMzMzMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzREREMzMzREREREREREREREREREREREREVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVREREREREREREMzMzMzMzMzMzMzMzIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzVVVVMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiERERIiIiIiIiERERERERERERIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzREREMzMzMzMzMzMzREREMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzREREMzMzREREREREREREREREREREVVVVREREREREVVVVVVVVd3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVREREMzMzREREREREREREREREREREREREREREREREMzMzREREREREREREREREREREVVVVZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREZmZmZmZmd3d3iIiId3d3d3d3d3d3ZmZmZmZmZmZmZmZmVVVVREREREREMzMzMzMzREREREREVVVVREREVVVVREREREREREREVVVVREREREREVVVVVVVVVVVVVVVVREREMzMzREREMzMzREREREREVVVVREREVVVVREREREREREREVVVVVVVVVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVZmZmZmZmd3d3ZmZmZmZmZmZmZmZmVVVVREREVVVVVVVVREREREREREREMzMzMzMzMzMzMzMzREREVVVVVVVVVVVVVVVVVVVVREREREREREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREMzMzREREREREVVVVVVVVZmZmd3d3ZmZmVVVVREREREREREREMzMzREREREREREREVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmVVVVREREREREREREREREMzMzMzMzMzMzMzMzREREREREREREREREREREREREVVVVVVVVZmZmVVVVREREMzMzMzMzMzMzREREMzMzMzMzMzMzREREMzMzMzMzMzMzREREVVVVVVVVVVVVVVVVZmZmVVVVVVVVREREMzMzREREREREMzMzREREREREMzMzREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVREREMzMzMzMzMzMzREREMzMzMzMzIiIiMzMzREREMzMzREREREREREREREREVVVVVVVVREREVVVVVVVVVVVVREREREREMzMzMzMzMzMzREREMzMzMzMzMzMzREREREREREREREREREREVVVVREREVVVVVVVVVVVVREREREREREREMzMzMzMzREREMzMzREREREREREREREREVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmd3d3d3d3VVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmREREREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3ZmZmZmZmVVVVVVVVVVVVREREVVVVVVVVZmZmd3d3iIiId3d3ZmZmVVVVREREVVVVVVVVVVVVZmZmZmZmd3d3d3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVd3d3d3d3d3d3d3d3ZmZmVVVVZmZmZmZmZmZmZmZmVVVVVVVVREREREREVVVVREREVVVVVVVVVVVVVVVVREREVVVVVVVVREREVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVZmZmZmZmVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3iIiIiIiIiIiImZmZiIiId3d3iIiImZmZu7u7u7u7u7u7zMzMzMzM3d3d7u7u////////////////////////////////////////////7u7u////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////93d3czMzN3d3e7u7szMzJmZmZmZmaqqqqqqqoiIiIiIiJmZmZmZmZmZmaqqqqqqqqqqqqqqqpmZmZmZmZmZmZmZmZmZmZmZmXd3d3d3d2ZmZmZmZmZmZnd3d4iIiJmZmaqqqqqqqru7u7u7u7u7u8zMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzLu7u7u7u7u7u7u7u6qqqpmZmYiIiIiIiIiIiHd3d2ZmZmZmZlVVVVVVVURERERERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzM0RERERERERERERERERERERERERERERERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVURERERERDMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERCIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERESIiIhERERERERERERERERERERERERERERERESIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERERERDMzM0RERERERERERERERERERERERERERDMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMyIiIjMzMzMzMyIiIiIiIiIiIjMzMzMzMzMzM0RERERERERERERERFVVVURERFVVVURERFVVVURERFVVVURERFVVVWZmZmZmZlVVVVVVVURERDMzM0RERERERERERERERERERDMzM0RERERERERERERERERERERERERERERERERERERERFVVVVVVVWZmZmZmZnd3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d3d3d3d3d2ZmZlVVVURERERERFVVVWZmZnd3d1VVVURERFVVVURERFVVVVVVVURERERERFVVVXd3d3d3d4iIiHd3d2ZmZnd3d2ZmZmZmZnd3d3d3d2ZmZlVVVURERERERDMzM0RERERERERERFVVVURERFVVVURERERERERERERERFVVVVVVVWZmZlVVVVVVVURERERERDMzM0RERDMzM0RERERERERERFVVVURERFVVVURERFVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVVVVVURERERERDMzMzMzM0RERDMzM0RERERERERERFVVVURERERERERERFVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZkRERFVVVURERERERERERERERERERERERERERERERDMzM0RERERERERERFVVVVVVVWZmZlVVVVVVVURERFVVVVVVVURERFVVVVVVVURERFVVVVVVVURERERERERERERERDMzM0RERFVVVVVVVWZmZmZmZnd3d1VVVURERERERERERERERDMzMzMzM0RERFVVVVVVVWZmZmZmZlVVVURERFVVVVVVVWZmZmZmZmZmZkRERERERERERDMzM0RERDMzMzMzM0RERERERERERERERERERERERERERFVVVVVVVWZmZlVVVURERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERERERFVVVVVVVVVVVVVVVWZmZlVVVVVVVURERERERERERERERERERERERDMzM0RERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVURERDMzM0RERDMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzM0RERERERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVURERDMzM0RERDMzMzMzMzMzMzMzM0RERERERERERERERERERERERERERERERFVVVURERFVVVURERERERDMzM0RERDMzM0RERDMzM0RERERERERERERERFVVVVVVVVVVVWZmZlVVVVVVVVVVVURERFVVVVVVVVVVVVVVVURERFVVVVVVVXd3d3d3d3d3d2ZmZlVVVURERFVVVURERGZmZmZmZmZmZnd3d2ZmZmZmZnd3d2ZmZlVVVURERFVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d1VVVVVVVWZmZlVVVVVVVWZmZmZmZnd3d3d3d2ZmZlVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZlVVVVVVVVVVVURERFVVVWZmZnd3d4iIiHd3d1VVVVVVVVVVVXd3d2ZmZmZmZlVVVVVVVURERERERERERERERFVVVVVVVVVVVURERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERFVVVVVVVWZmZmZmZmZmZmZmZlVVVWZmZmZmZlVVVWZmZnd3d2ZmZnd3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiJmZmZmZmbu7u8zMzMzMzN3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7MzMzMzMzu7u7d3d27u7uqqqqqqqqqqqqIiIiIiIiZmZmqqqq7u7uqqqqqqqqqqqq7u7u7u7u7u7u7u7u7u7u7u7uqqqqqqqqZmZmIiIh3d3eIiIh3d3d3d3d3d3eIiIiIiIiZmZmIiIiZmZmqqqq7u7u7u7u7u7vMzMzMzMy7u7uqqqqqqqqZmZmZmZmIiIh3d3d3d3dmZmZVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZVVVVERERERERERERERERERERVVVVVVVVVVVVVVVVmZmZVVVVmZmZVVVVmZmZVVVVERERVVVVEREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIREREREREiIiIREREiIiIREREiIiIiIiIREREiIiIREREiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNEREQzMzNEREQzMzNEREREREQzMzNEREREREQzMzNEREREREQzMzNEREREREQzMzNEREQzMzMzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzNEREREREQzMzNERERVVVVVVVVVVVVERERERERERERVVVVVVVVVVVVERERmZmZmZmZVVVVEREQzMzMzMzMiIiIzMzMzMzMzMzNERERERERERERERERVVVVERERERERERERVVVVERERERERVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZVVVVmZmZmZmZVVVWIiIh3d3dmZmZmZmZERERERERERERERERVVVVmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVVVVV3d3d3d3d3d3dmZmZVVVVmZmZmZmZmZmZ3d3eIiIh3d3dVVVVEREREREREREREREQzMzNERERERERERERVVVVERERERERERERERERERERVVVVmZmZVVVVEREREREREREREREQzMzMzMzNERERERERERERVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVmZmZVVVVmZmZmZmZVVVVEREREREREREQzMzNERERERERVVVVmZmZVVVVVVVVVVVVERERVVVVERERVVVVmZmZVVVVmZmZmZmZmZmZmZmZVVVVERERERERERERVVVVEREQzMzNERERERERERERERERERERERERERERERERVVVVVVVVmZmZmZmZVVVVVVVVmZmZmZmZVVVVEREREREREREREREREREREREREREQzMzNERERERERERERVVVVVVVV3d3d3d3dmZmZVVVVEREREREREREQzMzNERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVEREREREREREREREREREQzMzNERERERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVEREQzMzMzMzNEREQzMzMzMzMzMzMzMzNERERERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVERERERERERERERERERERERERERERERERVVVVERERVVVVERERVVVVmZmZmZmZERERVVVVVVVVVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNERERVVVVERERVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVEREQzMzNEREQzMzMzMzNEREREREQzMzNERERERERERERERERERERVVVVVVVVVVVVVVVVERERERERERERERERERERERERERERERERERERERERERERVVVVVVVVmZmZmZmZVVVVVVVVERERVVVVERERVVVVVVVVVVVVERERVVVVVVVV3d3d3d3dmZmZVVVVVVVVERERERERVVVVVVVVmZmZ3d3dmZmZmZmZmZmZmZmZ3d3dmZmZVVVVVVVVVVVVERERVVVVmZmZmZmZmZmZ3d3dmZmZmZmZmZmZVVVVmZmZmZmZVVVVmZmZ3d3d3d3dmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZ3d3dmZmZVVVVVVVVmZmZmZmZ3d3d3d3d3d3dmZmZVVVVVVVVmZmZmZmZmZmZVVVVERERERERVVVVVVVVVVVVERERmZmZmZmZVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVERERERERVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3eIiIh3d3d3d3d3d3d3d3eIiIiZmZmZmZmZmZm7u7u7u7vMzMzu7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////3d3dzMzM3d3d3d3dzMzMqqqqu7u7zMzMqqqqiIiIiIiImZmZqqqqqqqqiIiIiIiImZmZmZmZu7u7zMzMzMzMu7u7u7u7zMzMu7u7qqqqu7u7qqqqmZmZmZmZiIiImZmZiIiIiIiIiIiIiIiImZmZqqqqqqqqqqqqqqqqqqqqmZmZiIiIiIiIiIiIiIiId3d3d3d3ZmZmZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiImZmZiIiImZmZmZmZiIiImZmZiIiIiIiImZmZmZmZmZmZmZmZiIiId3d3d3d3ZmZmZmZmZmZmZmZmd3d3ZmZmVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVREREREREMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiMzMzMzMzIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiMzMzREREREREREREMzMzREREREREMzMzMzMzREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREREREMzMzREREVVVVREREREREREREREREREREREREREREVVVVMzMzREREVVVVREREMzMzMzMzMzMzMzMzREREMzMzREREREREREREREREREREVVVVREREREREREREREREVVVVREREREREREREREREREREREREMzMzREREREREREREREREREREVVVVZmZmd3d3ZmZmVVVVVVVVREREREREVVVVREREZmZmZmZmZmZmZmZmVVVVZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVZmZmd3d3iIiId3d3VVVVREREREREREREREREREREMzMzREREREREVVVVVVVVREREREREREREREREZmZmd3d3VVVVREREVVVVREREREREREREREREREREREREREREVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVREREREREMzMzREREREREREREZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVREREVVVVZmZmVVVVZmZmZmZmVVVVVVVVVVVVREREREREREREREREREREMzMzREREREREREREVVVVREREREREVVVVREREVVVVVVVVZmZmZmZmZmZmd3d3ZmZmVVVVREREREREMzMzMzMzMzMzMzMzREREREREREREREREREREVVVVZmZmiIiId3d3ZmZmVVVVREREREREMzMzREREREREREREREREREREVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmd3d3VVVVVVVVREREREREREREREREREREREREREREREREREREREREREREREREVVVVVVVVZmZmZmZmVVVVREREREREREREREREMzMzREREMzMzMzMzREREREREREREREREVVVVVVVVZmZmVVVVVVVVZmZmZmZmVVVVVVVVREREREREREREVVVVREREVVVVVVVVREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmVVVVREREREREMzMzMzMzREREMzMzREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREREREVVVVVVVVZmZmVVVVVVVVVVVVd3d3ZmZmVVVVVVVVREREVVVVREREVVVVVVVVREREVVVVVVVVZmZmZmZmZmZmZmZmVVVVVVVVREREREREVVVVVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3ZmZmVVVVVVVVZmZmZmZmVVVVZmZmd3d3d3d3ZmZmREREREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVZmZmREREVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmd3d3d3d3iIiIiIiIiIiIiIiImZmZmZmZqqqqu7u7u7u73d3d7u7u////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7szMzMzMzLu7u6qqqpmZmbu7u8zMzIiIiHd3d3d3d5mZmYiIiGZmZmZmZlVVVWZmZnd3d4iIiIiIiJmZmZmZmaqqqqqqqpmZmZmZmaqqqqqqqqqqqqqqqqqqqpmZmZmZmZmZmYiIiJmZmYiIiIiIiHd3d3d3d3d3d4iIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiJmZmZmZmZmZmZmZmaqqqqqqqru7u7u7u7u7u8zMzLu7u6qqqru7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqpmZmYiIiIiIiHd3d3d3d4iIiHd3d3d3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVURERERERERERDMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMyIiIiIiIhERESIiIhERESIiIhERESIiIiIiIiIiIhERESIiIiIiIhERESIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMyIiIiIiIjMzM0RERCIiIiIiIjMzMzMzMzMzMzMzM0RERDMzM1VVVVVVVVVVVTMzMzMzM0RERDMzM0RERDMzMzMzM0RERDMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMyIiIjMzMyIiIiIiIhERERERESIiIhERERERERERERERERERESIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERDMzM0RERDMzM0RERDMzM0RERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERFVVVURERERERERERERERDMzMzMzM0RERERERERERERERERERERERDMzM0RERDMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMzMzM0RERFVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVXd3d2ZmZlVVVURERERERFVVVVVVVVVVVXd3d2ZmZnd3d2ZmZlVVVURERERERERERERERERERERERFVVVURERERERERERERERERERFVVVWZmZoiIiGZmZkRERERERERERERERERERERERERERERERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVWZmZmZmZlVVVTMzM0RERERERFVVVVVVVVVVVURERERERERERERERFVVVURERFVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVURERERERERERERERDMzMzMzM0RERERERERERERERERERFVVVVVVVURERFVVVVVVVVVVVVVVVVVVVXd3d4iIiGZmZlVVVURERERERERERERERERERERERERERERERERERFVVVVVVVWZmZoiIiHd3d2ZmZmZmZlVVVURERERERFVVVURERERERERERERERERERERERFVVVVVVVWZmZmZmZmZmZnd3d3d3d3d3d2ZmZlVVVURERFVVVVVVVVVVVURERERERERERERERERERFVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVURERDMzM0RERERERDMzMzMzM0RERDMzM0RERERERERERFVVVVVVVVVVVWZmZmZmZnd3d2ZmZnd3d2ZmZlVVVVVVVURERFVVVURERERERFVVVURERFVVVURERFVVVURERFVVVURERFVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVURERERERERERERERDMzM0RERDMzM0RERERERERERERERFVVVVVVVURERFVVVVVVVVVVVVVVVWZmZmZmZnd3d2ZmZlVVVURERERERERERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVURERFVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZlVVVVVVVURERFVVVURERFVVVVVVVWZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZnd3d3d3d2ZmZmZmZmZmZlVVVWZmZnd3d4iIiGZmZmZmZmZmZlVVVVVVVXd3d3d3d3d3d3d3d4iIiGZmZlVVVVVVVVVVVURERFVVVVVVVVVVVWZmZlVVVURERERERFVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVWZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d5mZmZmZmaqqqqqqqru7u8zMzN3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7MzMy7u7uZmZmZmZmZmZmqqqqqqqqIiIhmZmZmZmZ3d3d3d3dmZmZmZmZmZmZVVVVmZmZ3d3dmZmaIiIiZmZmqqqqIiIh3d3d3d3eIiIh3d3d3d3d3d3d3d3eIiIh3d3eIiIiZmZmZmZmIiIiIiIiIiIiZmZmZmZmZmZmZmZmZmZmZmZmqqqqqqqq7u7uqqqqqqqq7u7uqqqq7u7u7u7u7u7u7u7u7u7u7u7uqqqqqqqqqqqq7u7u7u7uqqqq7u7u7u7u7u7uqqqqqqqqZmZmZmZmZmZmIiIiIiIiIiIhmZmZVVVVmZmZVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIzMzMiIiIiIiIiIiIiIiIREREiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzNERERERERVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIREREREREiIiIREREREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREQzMzNEREQzMzNEREREREREREQzMzNEREQzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzNERERERERVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERVVVVVVVVVVVVmZmZ3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZVVVVVVVVmZmZmZmZmZmZVVVVERERERERERERVVVVVVVVmZmZ3d3dmZmZVVVVERERERERERERERERVVVVERERVVVVERERERERVVVVERERERERVVVWIiIiZmZl3d3dVVVVERERERERERERERERVVVVERERVVVVVVVVVVVVVVVVVVVVERERERERERERVVVVmZmZmZmZmZmZmZmZmZmZ3d3dVVVVERERVVVVVVVVERERERERERERERERERERERERERERERERERERERERmZmZ3d3dmZmZmZmZVVVVmZmZVVVVVVVVEREREREREREREREREREQzMzMzMzNEREQzMzNERERERERVVVVERERVVVVVVVVmZmZmZmZmZmZVVVV3d3d3d3dVVVVVVVVERERERERERERERERERERERERERERERERERERVVVVVVVV3d3d3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERERERERERERERERERERERERERVVVVmZmZmZmZmZmZ3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERERERERERERERVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVERERERERERERVVVVERERERERERERERERERERERERVVVVERERERERmZmZmZmZmZmZ3d3dmZmZ3d3d3d3dVVVVVVVVERERVVVVERERVVVVERERERERERERERERVVVVERERVVVVVVVVVVVVmZmZVVVVmZmZmZmZ3d3dmZmZVVVVVVVVEREREREREREREREREREREREQzMzNERERERERVVVVVVVVVVVVVVVVVVVVERERERERVVVVVVVVVVVVmZmZmZmZVVVVVVVVERERVVVVERERERERERERVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3dmZmZVVVVVVVVmZmZmZmZmZmZmZmZ3d3eIiIh3d3dVVVVVVVVVVVVERERERERVVVVVVVVmZmZmZmZVVVVERERERERERERVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZVVVVmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZVVVVmZmZVVVVVVVVmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZmZmZ3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3eIiIiZmZmqqqrMzMzMzMzd3d3d3d3u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////3d3du7u7mZmZmZmZmZmZqqqqmZmZd3d3ZmZmZmZmd3d3d3d3ZmZmVVVVVVVVZmZmd3d3d3d3mZmZmZmZqqqqmZmZd3d3d3d3d3d3ZmZmZmZmd3d3iIiId3d3d3d3iIiImZmZmZmZmZmZmZmZu7u7u7u7qqqqu7u7u7u7qqqqu7u7u7u7qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqu7u7qqqqmZmZqqqqqqqqqqqqu7u7zMzMzMzMzMzMzMzMzMzMzMzMu7u7u7u7u7u7qqqqmZmZiIiIZmZmVVVVREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREVVVVREREREREMzMzMzMzREREREREMzMzMzMzMzMzREREMzMzIiIiIiIiMzMzMzMzMzMzIiIiIiIiMzMzIiIiERERERERERERERERERERERERIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzREREREREREREREREREREMzMzREREREREREREMzMzREREMzMzIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzREREMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREMzMzREREREREREREVVVVZmZmZmZmVVVVd3d3d3d3d3d3iIiId3d3d3d3VVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVREREVVVVREREVVVVVVVVZmZmZmZmZmZmVVVVVVVVREREREREREREREREVVVVREREREREREREREREREREREREVVVVd3d3mZmZZmZmREREREREVVVVVVVVREREREREVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmd3d3d3d3ZmZmZmZmZmZmVVVVREREREREREREREREMzMzREREREREREREREREMzMzREREVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVREREREREREREREREREREREREREREMzMzREREREREREREREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3d3d3VVVVVVVVREREREREREREREREREREREREREREVVVVVVVVVVVVZmZmd3d3d3d3ZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVREREVVVVVVVVVVVVREREVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3ZmZmZmZmREREREREVVVVVVVVREREVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVZmZmd3d3ZmZmZmZmZmZmZmZmZmZmVVVVREREREREREREVVVVREREREREREREREREVVVVREREVVVVVVVVZmZmVVVVZmZmVVVVVVVVZmZmZmZmZmZmVVVVVVVVREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVZmZmVVVVZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmVVVVVVVVZmZmVVVVVVVVZmZmZmZmVVVVZmZmVVVVZmZmZmZmZmZmZmZmd3d3ZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3ZmZmZmZmVVVVVVVVZmZmZmZmVVVVZmZmd3d3d3d3d3d3ZmZmVVVVREREVVVVVVVVVVVVREREZmZmd3d3ZmZmZmZmREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmVVVVVVVVZmZmZmZmVVVVZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmVVVVZmZmZmZmZmZmd3d3ZmZmZmZmVVVVZmZmZmZmd3d3ZmZmZmZmZmZmVVVVVVVVVVVVZmZmZmZmVVVVZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmd3d3ZmZmZmZmd3d3ZmZmZmZmd3d3iIiImZmZqqqqmZmZmZmZmZmZu7u73d3d3d3d////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7t3d3czMzLu7u6qqqqqqqqqqqru7u6qqqpmZmZmZmYiIiGZmZmZmZmZmZmZmZmZmZnd3d5mZmZmZmZmZmYiIiHd3d2ZmZmZmZmZmZnd3d4iIiHd3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d3d3d4iIiJmZmYiIiJmZmaqqqpmZmZmZmZmZmZmZmZmZmaqqqqqqqqqqqqqqqqqqqqqqqqqqqru7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqqqqqpmZmYiIiHd3d2ZmZkRERERERDMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIiIiAP//AAAiIiIiIiIiIiIiERERIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREREREREREREREMzMzREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzIiIiIiIiIiIiMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzREREMzMzREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREREREMzMzREREREREREREREREREREREREVVVVREREVVVVVVVVZmZmZmZmd3d3d3d3iIiIiIiId3d3VVVVVVVVVVVVZmZmVVVVd3d3d3d3iIiIZmZmVVVVZmZmZmZmZmZmZmZmZmZmVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmVVVVREREREREREREVVVVVVVVREREREREREREVVVVVVVVVVVVVVVVZmZmiIiId3d3VVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3VVVVREREREREREREREREREREREREMzMzREREREREREREVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREVVVVREREREREREREREREREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3ZmZmVVVVREREREREREREREREREREREREREREREREVVVVZmZmiIiId3d3ZmZmZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVREREREREREREVVVVZmZmd3d3d3d3ZmZmVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmVVVVVVVVREREVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVREREVVVVZmZmZmZmVVVVVVVVREREVVVVREREVVVVVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmVVVVREREVVVVVVVVZmZmZmZmd3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVZmZmVVVVVVVVREREREREMzMzREREREREREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREVVVVVVVVREREVVVVVVVVREREVVVVZmZmVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVZmZmZmZmVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmd3d3ZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmd3d3d3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVZmZmd3d3ZmZmZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmd3d3d3d3ZmZmZmZmVVVVZmZmd3d3d3d3ZmZmZmZmZmZmVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmd3d3d3d3d3d3d3d3d3d3iIiIiIiImZmZqqqqqqqqqqqqu7u7zMzM3d3d7u7u////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////+7u7u7u7t3d3d3d3czMzN3d3bu7u5mZmXd3d4iIiHd3d4iIiJmZmXd3d3d3d4iIiJmZmZmZmYiIiIiIiGZmZmZmZmZmZnd3d2ZmZmZmZlVVVXd3d3d3d3d3d2ZmZlVVVVVVVVVVVVVVVVVVVWZmZoiIiJmZmaqqqqqqqqqqqqqqqqqqqqqqqpmZmZmZmZmZmZmZmZmZmYiIiIiIiJmZmYiIiHd3d3d3d2ZmZnd3d2ZmZnd3d2ZmZlVVVVVVVURERERERDMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMyIiIjMzMyIiIiIiIjMzMyIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzM0RERDMzMzMzM0RERDMzMzMzM0RERDMzM0RERDMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzM0RERDMzM0RERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzMzMzMzMzMzMzMyIiIiIiIiIiIhERESIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMyIiIjMzMyIiIhERERERESIiIjMzM0RERERERERERDMzM0RERERERERERERERERERERERDMzM0RERERERERERERERERERERERFVVVURERDMzMzMzM0RERERERFVVVURERERERERERERERCIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzM0RERERERERERERERERERERERERERERERERERDMzM0RERERERDMzMzMzMzMzMzMzMzMzM0RERERERERERERERERERERERERERERERERERERERERERFVVVURERERERERERERERFVVVURERFVVVVVVVVVVVVVVVURERFVVVWZmZmZmZnd3d3d3d1VVVVVVVVVVVWZmZmZmZmZmZnd3d4iIiFVVVVVVVVVVVVVVVVVVVXd3d3d3d1VVVVVVVVVVVVVVVVVVVURERFVVVWZmZnd3d1VVVVVVVVVVVVVVVURERERERFVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d3d3d2ZmZlVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVWZmZmZmZnd3d4iIiHd3d4iIiHd3d4iIiHd3d2ZmZmZmZlVVVURERERERDMzM0RERERERERERFVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVVVVVVVVVURERFVVVURERERERFVVVURERERERERERFVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZlVVVURERERERFVVVURERERERFVVVVVVVVVVVWZmZnd3d3d3d1VVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d1VVVVVVVURERERERERERFVVVVVVVWZmZmZmZlVVVVVVVVVVVWZmZmZmZmZmZnd3d2ZmZnd3d2ZmZmZmZmZmZlVVVWZmZoiIiHd3d2ZmZlVVVURERERERFVVVURERFVVVVVVVURERFVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVURERFVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVURERFVVVVVVVVVVVWZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZlVVVWZmZlVVVVVVVVVVVVVVVURERERERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVURERERERFVVVURERFVVVVVVVURERFVVVURERFVVVVVVVVVVVWZmZlVVVURERFVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVWZmZlVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZnd3d2ZmZnd3d4iIiHd3d2ZmZmZmZlVVVVVVVWZmZlVVVVVVVWZmZmZmZnd3d3d3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVURERGZmZnd3d3d3d3d3d2ZmZmZmZlVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVURERFVVVVVVVWZmZnd3d2ZmZmZmZlVVVVVVVWZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZnd3d3d3d2ZmZnd3d4iIiIiIiIiIiHd3d3d3d4iIiJmZmaqqqru7u7u7u7u7u7u7u8zMzO7u7u7u7v///////////////////////////////////////////////////////////////////////+7u7v///////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3MzMyqqqqIiIiIiIiIiIh3d3eIiIh3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3d3d3dmZmZmZmZmZmZmZmZmZmaIiIh3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmaIiIiZmZmIiIiIiIiIiIh3d3dmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzNEREREREQzMzMzMzMzMzMzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzNEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNEREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMiIiIiIiIiIiIREREiIiIREREREREiIiIiIiIiIiIzMzMzMzNEREQzMzMzMzMzMzMiIiIiIiIREREiIiIiIiIiIiIiIiIzMzNERERVVVVERERERERVVVVEREREREREREQzMzNEREQzMzNERERVVVVVVVVERERERERERERVVVVEREREREQzMzMzMzNEREREREQzMzMiIiIzMzMiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzNERERERERVVVVVVVVVVVVVVVVVVVVEREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERVVVVEREREREREREREREREREREREQzMzNERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERVVVVVVVVVVVV3d3dmZmZmZmZVVVVVVVVmZmZmZmZVVVV3d3dmZmZVVVVERERVVVVVVVVVVVVmZmZ3d3dmZmZVVVVVVVVERERVVVVVVVVVVVVmZmZmZmZ3d3dmZmZVVVVERERVVVVERERVVVVVVVVmZmZmZmZmZmZVVVV3d3d3d3d3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVV3d3eIiIh3d3d3d3d3d3eIiIiIiIh3d3dmZmZmZmZmZmZVVVVERERERERERERERERERERVVVVVVVVmZmZmZmZmZmZmZmZ3d3dmZmZVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVmZmZ3d3d3d3dmZmZmZmZmZmZVVVVmZmZVVVVmZmZVVVVmZmZmZmZVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZVVVVmZmZVVVVmZmZVVVVmZmZ3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZVVVVVVVVVVVVmZmZ3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZ3d3dmZmZmZmZVVVVVVVVERERERERVVVVVVVVERERERERERERERERVVVVERERVVVVERERVVVVVVVVVVVVmZmZmZmZVVVVERERERERERERERERVVVVERERVVVVERERERERVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZVVVVmZmZmZmZ3d3dmZmZmZmZmZmZmZmZ3d3d3d3dVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZ3d3eIiIh3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVERERmZmZ3d3d3d3dmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3dmZmZ3d3d3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIiqqqrMzMzMzMzd3d3d3d3u7u7u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3dzMzMqqqqiIiId3d3ZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmVVVVREREREREREREREREMzMzMzMzREREREREMzMzREREREREREREREREMzMzMzMzREREREREREREREREMzMzMzMzMzMzREREREREREREREREREREREREREREMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzREREMzMzREREREREREREREREMzMzMzMzREREREREMzMzMzMzMzMzMzMzIiIiERERIiIiERERIiIiIiIiERERERERIiIiIiIiIiIiIiIiERERIiIiERERIiIiIiIiIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiMzMzREREVVVVREREREREREREVVVVVVVVMzMzMzMzREREMzMzMzMzREREREREMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzIiIiIiIiIiIiERERIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzREREREREREREREREVVVVVVVVREREVVVVREREREREMzMzMzMzMzMzMzMzMzMzREREREREMzMzREREREREREREREREREREREREMzMzREREMzMzMzMzREREMzMzMzMzREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVd3d3ZmZmd3d3VVVVVVVVVVVVZmZmVVVVd3d3d3d3iIiIZmZmZmZmVVVVZmZmVVVVVVVVZmZmZmZmVVVVVVVVd3d3ZmZmd3d3iIiIZmZmd3d3d3d3ZmZmZmZmVVVVVVVVVVVVZmZmVVVVVVVVVVVVZmZmVVVVVVVVZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmVVVVVVVVREREVVVVREREVVVVVVVVVVVVZmZmd3d3d3d3d3d3ZmZmZmZmVVVVVVVVREREVVVVREREVVVVZmZmZmZmZmZmZmZmVVVVVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmZmZmVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVREREREREREREZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3ZmZmZmZmd3d3d3d3d3d3d3d3ZmZmZmZmVVVVVVVVZmZmVVVVVVVVZmZmVVVVZmZmVVVVVVVVZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVREREVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVREREVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVREREZmZmZmZmZmZmd3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREVVVVZmZmZmZmZmZmZmZmVVVVREREREREREREREREVVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmVVVVZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmVVVVd3d3ZmZmZmZmVVVVZmZmZmZmd3d3ZmZmZmZmZmZmVVVVVVVVVVVVREREVVVVZmZmZmZmd3d3d3d3d3d3d3d3ZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmd3d3d3d3ZmZmVVVVVVVVZmZmZmZmZmZmd3d3VVVVZmZmVVVVVVVVVVVVVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmZmZmd3d3ZmZmZmZmZmZmd3d3d3d3iIiIiIiId3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiIqqqqu7u73d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7t3d3czMzJmZmYiIiHd3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERERERERERERERFVVVURERERERFVVVVVVVWZmZmZmZlVVVXd3d3d3d3d3d3d3d4iIiJmZmZmZmZmZmZmZmZmZmaqqqpmZmZmZmaqqqpmZmZmZmZmZmZmZmYiIiIiIiIiIiGZmZmZmZlVVVVVVVVVVVTMzM0RERERERERERDMzM0RERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIhERESIiIhERESIiIiIiIiIiIhERERERERERERERERERESIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMyIiIjMzM0RERERERDMzM0RERDMzMzMzM0RERERERFVVVVVVVTMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERERERDMzM0RERERERDMzMzMzMzMzM0RERERERDMzMzMzM0RERERERERERDMzM0RERERERERERERERDMzM0RERERERERERERERDMzM0RERDMzM0RERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVXd3d4iIiIiIiHd3d2ZmZmZmZnd3d3d3d3d3d3d3d1VVVVVVVURERERERGZmZnd3d2ZmZmZmZnd3d2ZmZnd3d3d3d4iIiIiIiGZmZlVVVWZmZlVVVWZmZmZmZnd3d3d3d2ZmZlVVVWZmZnd3d3d3d3d3d4iIiHd3d2ZmZnd3d3d3d3d3d2ZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVWZmZmZmZnd3d3d3d4iIiHd3d2ZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d3d3d3d3d2ZmZlVVVURERFVVVURERFVVVVVVVWZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZnd3d2ZmZlVVVURERERERFVVVWZmZlVVVURERFVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZlVVVVVVVVVVVURERERERFVVVURERFVVVWZmZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZlVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d2ZmZnd3d2ZmZmZmZlVVVVVVVVVVVWZmZlVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVWZmZnd3d2ZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVURERFVVVURERFVVVWZmZnd3d2ZmZnd3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVURERFVVVURERERERFVVVVVVVURERERERFVVVVVVVWZmZmZmZmZmZnd3d2ZmZlVVVURERERERERERFVVVURERFVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVWZmZmZmZnd3d3d3d4iIiJmZmaqqqoiIiHd3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d1VVVVVVVVVVVWZmZmZmZnd3d3d3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZnd3d3d3d4iIiGZmZlVVVVVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVURERFVVVVVVVVVVVWZmZlVVVWZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVWZmZmZmZlVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d2ZmZmZmZnd3d3d3d3d3d4iIiHd3d3d3d3d3d4iIiJmZmZmZmZmZmYiIiIiIiHd3d5mZmaqqqqqqqpmZmaqqqru7u8zMzO7u7u7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////u7u7d3d2qqqqIiIh3d3d3d3d3d3dmZmZ3d3d3d3d3d3d3d3eIiIh3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZ3d3d3d3d3d3eIiIiZmZmZmZmZmZmqqqq7u7u7u7uqqqq7u7u7u7uqqqq7u7u7u7u7u7u7u7uqqqqqqqqqqqqIiIiIiIhmZmZmZmZVVVVERERVVVVERERERERERERERERVVVVERERERERERERVVVVERERERERERERVVVVEREREREQzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIREREiIiIREREREREiIiIREREiIiIREREREREiIiIiIiIREREiIiIREREiIiIiIiIzMzMiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNEREREREQzMzMiIiIREREiIiIREREREREREREiIiIiIiIzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzNERERVVVVEREREREREREQzMzNEREREREQzMzNEREREREQzMzMzMzMzMzNEREREREREREQzMzNEREREREQzMzMzMzNEREREREQzMzMzMzMzMzNEREREREREREREREREREREREREREREREREREQzMzNEREQzMzNEREQzMzNERERERERERERVVVVVVVVVVVVERERVVVVVVVVERERVVVVERERVVVVVVVWIiIiZmZmZmZmIiIh3d3d3d3eIiIh3d3d3d3d3d3d3d3dVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3eIiIiIiIhmZmaIiIh3d3dmZmZVVVVVVVVVVVVVVVVmZmZ3d3dmZmZVVVVmZmZmZmZ3d3dmZmaIiIh3d3dmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVmZmZVVVVmZmZmZmZ3d3eIiIhmZmZmZmZmZmZVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3d3d3eIiIh3d3eIiIh3d3eIiIh3d3dmZmZVVVVVVVVVVVVERERVVVVVVVVmZmZVVVVVVVVmZmZ3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3eIiIiIiIh3d3dmZmZERERVVVVVVVVERERERERVVVVERERVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZmZmZVVVVmZmZVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZVVVVmZmZmZmZmZmZmZmZ3d3dmZmZ3d3dVVVVVVVVVVVVmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3dmZmZ3d3d3d3dmZmZVVVVVVVVERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERERERVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERERERVVVVERERVVVVmZmaIiIi7u7uqqqqqqqp3d3d3d3dmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmaIiIh3d3dmZmZVVVVmZmZVVVVmZmZmZmaIiIh3d3d3d3dmZmZVVVVVVVVmZmZVVVVVVVVERERVVVVmZmZmZmZ3d3dmZmZmZmZVVVVmZmZVVVVmZmZVVVVmZmZmZmZVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZVVVVmZmZmZmZVVVVmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZVVVVmZmZVVVVmZmZmZmZmZmZ3d3d3d3dmZmZmZmZ3d3d3d3eIiIh3d3eIiIh3d3eIiIiIiIiqqqqZmZmZmZmZmZmZmZmZmZm7u7vMzMzd3d3d3d3MzMzd3d3u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////3d3dzMzMu7u7mZmZiIiId3d3d3d3d3d3d3d3iIiIiIiImZmZmZmZiIiIiIiImZmZmZmZmZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZmZmZqqqqqqqqu7u7qqqqu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7qqqqqqqqiIiId3d3ZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVZmZmREREREREREREVVVVREREMzMzMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiERERIiIiERERIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzREREMzMzREREMzMzREREMzMzREREREREMzMzMzMzMzMzIiIiIiIiIiIiMzMzIiIiMzMzMzMzIiIiIiIiIiIiIiIiERERIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREREREREREREREREREREREMzMzMzMzREREREREREREMzMzREREMzMzMzMzREREMzMzREREREREREREREREREREMzMzMzMzMzMzREREMzMzMzMzMzMzVVVVREREMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREVVVVVVVVVVVVVVVVREREVVVVREREREREREREZmZmZmZmmZmZiIiId3d3iIiId3d3d3d3iIiId3d3iIiId3d3d3d3ZmZmREREVVVVZmZmd3d3ZmZmd3d3d3d3iIiImZmZiIiId3d3d3d3d3d3d3d3ZmZmREREVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmd3d3ZmZmZmZmZmZmZmZmVVVVZmZmZmZmd3d3d3d3iIiId3d3ZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiIZmZmVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmZmZmd3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmd3d3ZmZmVVVVVVVVZmZmZmZmd3d3d3d3iIiIiIiId3d3ZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmd3d3d3d3VVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmREREVVVVVVVVZmZmVVVVZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmVVVVZmZmVVVVZmZmd3d3VVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmVVVVZmZmd3d3ZmZmd3d3ZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVREREVVVVREREVVVVVVVVREREVVVVVVVVREREREREREREREREMzMzMzMzREREMzMzREREREREREREVVVViIiIqqqqmZmZiIiId3d3d3d3ZmZmd3d3d3d3ZmZmd3d3ZmZmZmZmVVVVVVVVZmZmZmZmZmZmZmZmd3d3d3d3ZmZmZmZmmZmZiIiIZmZmVVVVZmZmZmZmZmZmd3d3iIiIiIiIZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVREREVVVVVVVVZmZmZmZmVVVVZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3iIiId3d3d3d3d3d3iIiImZmZmZmZiIiIiIiImZmZmZmZqqqqqqqqqqqqmZmZqqqqu7u7zMzM7u7u7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////+7u7u7u7t3d3d3d3bu7u5mZmXd3d2ZmZlVVVWZmZmZmZmZmZmZmZoiIiIiIiIiIiKqqqpmZmaqqqqqqqqqqqqqqqqqqqru7u6qqqru7u7u7u7u7u7u7u7u7u8zMzLu7u7u7u8zMzMzMzLu7u7u7u7u7u7u7u6qqqpmZmZmZmYiIiHd3d2ZmZnd3d2ZmZlVVVURERERERFVVVURERERERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMyIiIjMzMyIiIjMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMyIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMyIiIjMzMzMzMyIiIjMzMyIiIiIiIiIiIjMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIjMzMzMzMzMzMyIiIjMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERERERDMzM0RERDMzM0RERDMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIhERESIiIhERERERERERERERESIiIhERESIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIjMzMzMzMzMzM0RERDMzM0RERDMzMzMzM0RERERERERERERERDMzM0RERDMzMzMzM0RERERERERERERERDMzMzMzMzMzMzMzM0RERERERDMzMzMzMzMzMzMzMzMzM0RERERERERERDMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERERERFVVVVVVVVVVVURERERERERERERERERERERERFVVVXd3d4iIiGZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZnd3d3d3d2ZmZmZmZlVVVWZmZnd3d4iIiHd3d3d3d4iIiIiIiIiIiGZmZmZmZnd3d4iIiHd3d2ZmZlVVVVVVVWZmZmZmZnd3d2ZmZlVVVWZmZmZmZnd3d3d3d3d3d3d3d3d3d2ZmZmZmZmZmZnd3d3d3d3d3d4iIiHd3d3d3d3d3d2ZmZnd3d2ZmZmZmZmZmZmZmZnd3d4iIiIiIiHd3d3d3d2ZmZlVVVVVVVVVVVWZmZlVVVWZmZmZmZnd3d4iIiIiIiHd3d4iIiIiIiIiIiIiIiGZmZlVVVVVVVWZmZnd3d2ZmZmZmZnd3d3d3d3d3d3d3d3d3d2ZmZmZmZnd3d2ZmZmZmZnd3d3d3d1VVVVVVVVVVVWZmZmZmZlVVVWZmZnd3d3d3d3d3d2ZmZnd3d2ZmZnd3d3d3d3d3d3d3d4iIiHd3d2ZmZlVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVWZmZlVVVWZmZmZmZnd3d3d3d2ZmZnd3d2ZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZnd3d3d3d2ZmZnd3d2ZmZnd3d3d3d2ZmZlVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d2ZmZlVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVURERFVVVVVVVVVVVURERFVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVURERERERFVVVURERERERFVVVVVVVVVVVURERFVVVURERERERERERFVVVURERERERERERDMzM0RERERERDMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIkRERHd3d4iIiIiIiIiIiHd3d3d3d2ZmZnd3d2ZmZnd3d2ZmZmZmZmZmZlVVVVVVVYiIiHd3d2ZmZmZmZmZmZnd3d2ZmZmZmZnd3d1VVVWZmZmZmZmZmZnd3d3d3d4iIiIiIiGZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVURERFVVVVVVVURERFVVVURERFVVVURERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZnd3d4iIiIiIiJmZmYiIiIiIiIiIiJmZmZmZmZmZmZmZmZmZmaqqqqqqqszMzMzMzLu7u7u7u8zMzN3d3e7u7v///////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7MzMy7u7uIiIhmZmZVVVVVVVVVVVVVVVVmZmZ3d3dmZmaIiIiIiIiIiIiIiIiZmZmZmZmZmZmZmZmZmZmZmZmZmZmqqqqqqqqqqqqqqqq7u7u7u7u7u7u7u7uqqqqZmZmqqqqqqqqqqqqZmZmZmZmIiIh3d3dmZmZVVVVEREREREQzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMiIiIzMzMiIiIzMzMiIiIzMzMzMzMiIiIzMzMiIiIiIiIzMzMzMzMiIiIzMzMiIiIiIiIzMzMzMzMzMzMiIiIiIiIzMzMzMzMiIiIzMzMzMzMiIiIzMzMiIiIiIiIzMzMiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzNEREREREQzMzNEREQzMzMzMzNEREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIREREiIiIiIiIREREiIiIiIiIREREiIiIREREiIiIiIiIiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREQzMzMzMzNEREQzMzMzMzMzMzNERERERERERERVVVVVVVVEREREREQzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREREREREREREREREREREREQzMzNEREQzMzNEREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERERERERERERERVVVVVVVVVVVVVVVVEREREREQzMzNVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVEREREREQzMzNERERVVVVmZmZ3d3dmZmZ3d3d3d3dmZmZmZmZ3d3d3d3dmZmZ3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3d3d3d3d3dmZmZmZmZVVVVmZmZmZmZ3d3d3d3d3d3dmZmZmZmZmZmZ3d3d3d3d3d3eIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIiZmZmIiIiIiIiIiIh3d3dmZmZVVVVmZmZVVVVVVVVmZmZmZmZ3d3eIiIiZmZmZmZmZmZmIiIiIiIiIiIh3d3dmZmZVVVVVVVV3d3d3d3d3d3d3d3d3d3eIiIh3d3eZmZmIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3dmZmZmZmZmZmZVVVVmZmZmZmZ3d3d3d3eIiIh3d3d3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3eIiIh3d3dVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3eIiIh3d3d3d3dmZmZmZmZmZmZmZmZ3d3d3d3dmZmZ3d3dmZmZ3d3dmZmZ3d3d3d3dmZmZ3d3dmZmZ3d3d3d3d3d3dVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZVVVVVVVVmZmZmZmZmZmZmZmZ3d3d3d3dmZmZmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3dmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERERERERERVVVVERERERERVVVVERERERERERERERERERERERERERERVVVVEREREREREREREREQzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiJERERmZmZ3d3dVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVERERmZmaIiIh3d3dVVVVVVVVVVVVmZmZmZmZmZmZVVVVVVVVmZmZ3d3dmZmZmZmZ3d3d3d3d3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVERERERERVVVVVVVVmZmZVVVVERERERERERERVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3dmZmZ3d3eIiIh3d3d3d3d3d3d3d3eIiIiIiIiIiIiZmZmIiIiZmZmIiIiZmZmZmZmIiIiZmZmZmZmqqqqqqqq7u7vMzMzd3d3d3d3d3d3u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////7u7u////////////////////////////////////////7u7u7u7uu7u7mZmZd3d3ZmZmd3d3ZmZmZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmd3d3iIiId3d3mZmZmZmZmZmZmZmZiIiImZmZqqqqqqqqmZmZmZmZqqqqmZmZmZmZmZmZqqqqmZmZiIiId3d3ZmZmVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiIiIiIiIiMzMzMzMzIiIiMzMzIiIiMzMzMzMzIiIiMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzIiIiMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVREREREREMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiERERIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREMzMzREREREREREREMzMzREREREREVVVVVVVVVVVVVVVVVVVVREREREREMzMzREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREREREREREMzMzREREMzMzMzMzREREREREMzMzREREREREMzMzREREREREREREMzMzREREREREREREREREVVVVREREREREREREVVVVREREZmZmZmZmVVVVVVVVREREREREREREREREREREREREREREREREREREVVVVVVVVZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmVVVVZmZmd3d3d3d3d3d3ZmZmZmZmd3d3iIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmd3d3ZmZmiIiId3d3d3d3d3d3ZmZmd3d3d3d3d3d3iIiIiIiIiIiId3d3iIiIiIiId3d3iIiIiIiImZmZmZmZmZmZiIiId3d3ZmZmZmZmVVVVVVVVVVVVZmZmZmZmd3d3iIiIqqqqmZmZqqqqmZmZiIiIiIiIiIiIiIiId3d3ZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiImZmZmZmZmZmZmZmZiIiIiIiIiIiId3d3iIiIiIiIZmZmZmZmVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiId3d3iIiIiIiId3d3ZmZmVVVVZmZmVVVVVVVVZmZmZmZmVVVVZmZmd3d3d3d3d3d3iIiId3d3d3d3d3d3iIiIZmZmZmZmd3d3d3d3ZmZmd3d3iIiId3d3d3d3iIiId3d3d3d3ZmZmZmZmd3d3ZmZmd3d3d3d3ZmZmZmZmVVVVZmZmVVVVZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVZmZmVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVREREREREREREREREREREREREREREREREREREREREREREREREMzMzMzMzREREREREREREREREREREREREREREMzMzMzMzMzMzIiIiIiIiIiIiMzMzIiIiMzMzIiIiIiIiMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVREREMzMzMzMzMzMzMzMzREREREREREREREREMzMzMzMzREREZmZmVVVVREREREREREREVVVVVVVVZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREZmZmZmZmVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmiIiId3d3d3d3iIiId3d3d3d3d3d3mZmZiIiIiIiImZmZmZmZmZmZmZmZmZmZiIiIiIiImZmZiIiImZmZqqqqqqqqqqqqqqqqu7u7u7u73d3d3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////93d3bu7u5mZmYiIiIiIiJmZmZmZmZmZmYiIiIiIiHd3d2ZmZnd3d2ZmZmZmZmZmZnd3d4iIiIiIiIiIiIiIiIiIiIiIiJmZmZmZmZmZmYiIiIiIiJmZmYiIiIiIiIiIiIiIiHd3d2ZmZlVVVURERERERDMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzM0RERGZmZmZmZkRERDMzMzMzMyIiIiIiIiIiIhERESIiIhERESIiIhERESIiIiIiIjMzMyIiIjMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzM0RERDMzM0RERDMzMzMzM0RERERERDMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM0RERERERFVVVURERERERDMzM0RERDMzM0RERERERERERERERERERERERERERERERFVVVVVVVTMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzMzMzM0RERERERDMzM0RERERERERERDMzM0RERERERERERERERERERERERERERFVVVVVVVURERFVVVVVVVURERERERERERDMzMzMzM0RERERERFVVVVVVVVVVVURERFVVVVVVVVVVVWZmZmZmZoiIiIiIiIiIiIiIiHd3d3d3d1VVVWZmZnd3d3d3d4iIiHd3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiIiIiHd3d3d3d2ZmZmZmZmZmZoiIiJmZmZmZmXd3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiIiIiHd3d3d3d3d3d4iIiIiIiJmZmYiIiIiIiIiIiHd3d4iIiHd3d2ZmZmZmZmZmZmZmZmZmZnd3d4iIiKqqqpmZmZmZmYiIiIiIiHd3d3d3d4iIiHd3d2ZmZmZmZmZmZmZmZmZmZnd3d4iIiIiIiJmZmZmZmZmZmZmZmYiIiIiIiHd3d4iIiHd3d4iIiHd3d1VVVWZmZlVVVWZmZmZmZmZmZmZmZnd3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiIiIiHd3d2ZmZmZmZmZmZnd3d2ZmZmZmZnd3d3d3d3d3d3d3d4iIiIiIiHd3d3d3d4iIiHd3d4iIiHd3d2ZmZnd3d3d3d3d3d3d3d4iIiHd3d4iIiIiIiHd3d3d3d2ZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVURERGZmZlVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERDMzMzMzM0RERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMyIiIiIiIjMzMzMzMyIiIjMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzM0RERDMzM0RERERERDMzMzMzM0RERDMzMzMzM0RERERERERERDMzMzMzM0RERERERERERERERERERERERERERERERDMzM0RERERERFVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZlVVVURERERERFVVVVVVVVVVVWZmZlVVVWZmZmZmZlVVVVVVVURERERERFVVVVVVVVVVVURERFVVVVVVVURERFVVVVVVVVVVVVVVVURERFVVVVVVVWZmZlVVVVVVVWZmZmZmZmZmZmZmZmZmZnd3d4iIiJmZmYiIiJmZmYiIiIiIiJmZmaqqqpmZmaqqqpmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmaqqqru7u8zMzMzMzN3d3d3d3d3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7MzMy7u7uqqqqqqqqqqqq7u7u7u7u7u7uZmZmZmZmZmZmqqqqZmZmZmZmIiIiIiIiIiIiIiIh3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZmIiIiIiIh3d3d3d3dmZmZmZmZmZmZ3d3dmZmZVVVVVVVVmZmZVVVVVVVVERERVVVVVVVVEREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERVVVVEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNEREQzMzNEREQzMzNEREREREREREQzMzNEREQzMzNEREQzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzNERER3d3dmZmZEREQzMzMiIiIiIiIiIiIiIiIREREiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMiIiIzMzMzMzNERERERERERERVVVVEREREREREREREREQzMzNEREREREREREREREREREREREREREQzMzNERERERERERERVVVVERERVVVVEREQzMzMzMzMzMzMiIiIzMzMzMzMzMzNEREQzMzNERERVVVVVVVVEREREREREREREREREREQzMzMzMzNEREQzMzMzMzMzMzNEREREREREREQzMzNEREREREQzMzNERERERERERERVVVVEREREREQzMzMzMzNEREQzMzNERERERERVVVVVVVVVVVVVVVVVVVVVVVVEREREREREREREREQzMzNERERERERVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVmZmZmZmZ3d3d3d3eZmZmZmZmZmZmIiIiIiIh3d3d3d3eIiIiIiIh3d3eIiIh3d3eIiIh3d3eIiIiIiIiIiIh3d3eIiIiIiIiIiIh3d3d3d3d3d3dmZmZ3d3d3d3eIiIh3d3eIiIiIiIiIiIiIiIh3d3d3d3d3d3eIiIh3d3d3d3eIiIh3d3d3d3d3d3eIiIiIiIh3d3eIiIh3d3eIiIiZmZmZmZmIiIh3d3d3d3d3d3d3d3d3d3d3d3eIiIiZmZmZmZmIiIiIiIh3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIiIiIiZmZmZmZmIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3dmZmZ3d3dmZmZ3d3eIiIh3d3d3d3eIiIiIiIiIiIh3d3d3d3d3d3d3d3eIiIiIiIh3d3dmZmZ3d3d3d3d3d3d3d3dmZmZ3d3eIiIiIiIh3d3d3d3dmZmaIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3dmZmZ3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZVVVVmZmZ3d3dmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZ3d3dmZmZmZmZVVVVVVVVmZmZmZmZmZmZmZmZVVVVmZmZVVVVVVVVmZmZVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVmZmZVVVVVVVVmZmZVVVVmZmZVVVVmZmZVVVVmZmZVVVVVVVVVVVVVVVVERERVVVVERERVVVVEREREREREREREREREREREREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMiIiIiIiIiIiIzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzNERERERERERERERERERERERERERERVVVVERERERERERERVVVVEREREREREREREREREREREREQzMzNEREQzMzNERERERERERERERERERERERERERERERERERERVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZVVVVVVVVVVVVERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVmZmZmZmZ3d3d3d3d3d3eIiIiIiIh3d3eIiIiZmZmZmZmZmZmZmZmZmZmqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqq7u7u7u7u7u7vMzMzd3d3d3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3du7u7u7u7u7u7u7u7u7u7u7u7zMzMzMzMzMzMzMzMzMzMu7u7qqqqqqqqu7u7qqqqqqqqqqqqqqqqqqqqqqqqqqqqu7u7qqqqu7u7qqqqu7u7qqqqqqqqqqqqqqqqqqqqqqqqqqqqmZmZmZmZiIiImZmZiIiId3d3iIiIiIiId3d3d3d3ZmZmVVVVREREMzMzMzMzMzMzREREMzMzREREREREMzMzMzMzREREREREREREREREREREVVVVVVVVREREREREMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzREREMzMzREREMzMzREREMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVd3d3d3d3REREMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREREREVVVVREREREREREREREREREREREREREREVVVVZmZmVVVVREREREREREREREREVVVVVVVVVVVVREREVVVVREREMzMzREREMzMzREREMzMzREREMzMzMzMzMzMzVVVVZmZmVVVVVVVVVVVVREREREREREREREREMzMzREREMzMzMzMzREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREREVVVVVVVVZmZmZmZmVVVVZmZmVVVVREREREREREREREREREREREREVVVVVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmd3d3iIiIiIiImZmZiIiIiIiIiIiIiIiIiIiIiIiImZmZiIiIiIiIiIiIiIiIiIiIiIiId3d3iIiIiIiIiIiId3d3iIiIiIiIiIiId3d3d3d3d3d3iIiIiIiIiIiId3d3d3d3iIiIiIiIiIiIiIiId3d3d3d3iIiIiIiIiIiIiIiIiIiId3d3iIiId3d3iIiIiIiIiIiIiIiImZmZqqqqmZmZmZmZiIiImZmZiIiId3d3d3d3d3d3iIiIiIiImZmZmZmZiIiId3d3d3d3iIiImZmZmZmZiIiImZmZiIiIiIiIiIiIiIiIiIiImZmZiIiIiIiId3d3iIiIiIiIiIiId3d3d3d3ZmZmd3d3iIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3iIiIiIiIiIiIiIiId3d3d3d3ZmZmd3d3d3d3d3d3iIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3iIiIiIiImZmZmZmZmZmZmZmZmZmZmZmZiIiImZmZiIiImZmZiIiId3d3d3d3d3d3d3d3d3d3iIiIiIiId3d3iIiId3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmd3d3d3d3VVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmREREVVVVREREVVVVREREREREREREREREREREREREREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzREREVVVVMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREVVVVVVVVVVVVREREVVVVREREVVVVVVVVVVVVREREVVVVVVVVREREMzMzREREREREREREREREREREVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREVVVVREREREREVVVVREREVVVVVVVVZmZmVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3iIiIiIiIiIiIiIiIiIiImZmZmZmZmZmZmZmZmZmZmZmZqqqqqqqqqqqqqqqqqqqqqqqqqqqqu7u7u7u7u7u7u7u7u7u7u7u7zMzM3d3d3d3d7u7u7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////+7u7t3d3czMzMzMzLu7u7u7u7u7u8zMzMzMzMzMzLu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u8zMzMzMzLu7u7u7u8zMzLu7u7u7u7u7u8zMzLu7u6qqqqqqqqqqqqqqqpmZmZmZmaqqqpmZmZmZmZmZmaqqqpmZmZmZmZmZmXd3d1VVVURERFVVVVVVVURERFVVVURERERERERERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzM0RERDMzM0RERDMzM0RERDMzM0RERDMzM0RERDMzMzMzMzMzM0RERERERDMzM0RERDMzM0RERDMzM0RERGZmZnd3d2ZmZkRERDMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzMzMzM0RERERERERERERERFVVVVVVVVVVVVVVVVVVVURERFVVVVVVVURERGZmZlVVVVVVVVVVVURERERERERERFVVVWZmZmZmZlVVVURERFVVVVVVVURERDMzMzMzMzMzMzMzMzMzMzMzM0RERERERERERFVVVWZmZmZmZlVVVWZmZlVVVURERERERERERERERDMzM0RERERERERERFVVVVVVVURERDMzM0RERERERERERERERFVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZkRERERERERERERERFVVVVVVVWZmZmZmZnd3d2ZmZmZmZmZmZmZmZlVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZoiIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiJmZmZmZmZmZmYiIiIiIiHd3d4iIiHd3d4iIiIiIiIiIiHd3d5mZmYiIiIiIiIiIiHd3d3d3d4iIiJmZmZmZmZmZmYiIiIiIiIiIiIiIiIiIiIiIiJmZmYiIiIiIiHd3d3d3d4iIiIiIiIiIiHd3d4iIiIiIiIiIiJmZmaqqqqqqqqqqqqqqqpmZmZmZmZmZmZmZmYiIiIiIiJmZmZmZmZmZmZmZmYiIiIiIiIiIiIiIiJmZmaqqqpmZmZmZmZmZmYiIiIiIiIiIiIiIiJmZmZmZmYiIiHd3d4iIiIiIiIiIiIiIiHd3d2ZmZnd3d4iIiHd3d4iIiIiIiIiIiHd3d3d3d3d3d4iIiHd3d4iIiHd3d4iIiIiIiHd3d2ZmZnd3d3d3d4iIiHd3d4iIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d3d3d4iIiIiIiIiIiHd3d4iIiJmZmZmZmZmZmaqqqqqqqqqqqru7u6qqqqqqqpmZmZmZmZmZmZmZmZmZmYiIiIiIiIiIiIiIiIiIiJmZmYiIiHd3d4iIiHd3d4iIiHd3d3d3d2ZmZnd3d3d3d3d3d3d3d2ZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVURERFVVVURERFVVVURERERERERERERERERERERERERERERERERERERERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIjMzMyIiIiIiIiIiIiIiIjMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzMyIiIjMzMyIiIjMzM0RERFVVVVVVVVVVVVVVVVVVVURERERERDMzMzMzM0RERERERFVVVURERERERERERERERDMzM0RERERERDMzMzMzMzMzMzMzM0RERERERERERERERERERERERERERFVVVURERFVVVVVVVVVVVVVVVVVVVVVVVVVVVURERERERFVVVURERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVURERERERFVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d2ZmZmZmZmZmZnd3d2ZmZmZmZnd3d3d3d4iIiIiIiIiIiJmZmYiIiJmZmZmZmaqqqpmZmZmZmaqqqqqqqqqqqru7u6qqqqqqqru7u8zMzMzMzN3d3d3d3d3d3d3d3e7u7u7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7d3d3MzMzMzMyqqqq7u7vMzMy7u7u7u7uqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqZmZmqqqqZmZmqqqqqqqqqqqq7u7uqqqqqqqq7u7u7u7u7u7uqqqqqqqqqqqqqqqqIiIh3d3dmZmZmZmZVVVVVVVVEREREREREREQzMzMzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIzMzMiIiIzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzMzMzNEREQzMzMzMzMzMzMzMzNEREREREQzMzNEREQzMzNEREREREREREREREREREQzMzMzMzNEREQzMzMzMzMzMzNERERVVVVVVVVVVVVVVVUzMzMiIiIiIiIzMzMiIiIiIiIzMzMzMzMzMzMzMzMiIiIzMzMzMzNEREQzMzNEREQzMzNEREQzMzMzMzNEREQzMzMzMzMzMzMzMzNERERERERERERVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZVVVVVVVVERERmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZERERERERERERERERERERVVVVERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVERERVVVVERERVVVVERERERERVVVVERERERERERERVVVVmZmZmZmZmZmZ3d3eIiIiIiIh3d3eIiIhmZmZmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZ3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3eIiIiIiIiZmZmZmZmIiIiIiIiIiIiIiIiZmZmIiIiIiIh3d3d3d3d3d3dmZmZ3d3d3d3d3d3eIiIiZmZmZmZmZmZmZmZmZmZmZmZmIiIiZmZmZmZmqqqqZmZmqqqqqqqqqqqqqqqqZmZmZmZmZmZmZmZmIiIh3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZmqqqqqqqqqqqqqqqqZmZmZmZmqqqqZmZmqqqqZmZmqqqqZmZmqqqqqqqqZmZmIiIiIiIiZmZmqqqqqqqqqqqqZmZmZmZmIiIiZmZmZmZmZmZmZmZmZmZmIiIiIiIiIiIiIiIiZmZl3d3d3d3d3d3eIiIiZmZmIiIiIiIiZmZmZmZmIiIiIiIiIiIiIiIh3d3d3d3eIiIiIiIiIiIh3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIiZmZmIiIiZmZmIiIiIiIh3d3eIiIiZmZmZmZmZmZmZmZmqqqq7u7u7u7u7u7u7u7u7u7u7u7u7u7vMzMy7u7uqqqqZmZmZmZmZmZmZmZmIiIiIiIiIiIiIiIiIiIh3d3eIiIh3d3d3d3d3d3dmZmZ3d3dmZmZmZmZmZmZ3d3d3d3dmZmZmZmZVVVVmZmZmZmZVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVEREREREREREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIzMzMzMzMzMzMzMzMiIiIzMzMiIiIiIiIiIiIzMzMzMzNEREQzMzMzMzMiIiIzMzMiIiIzMzMzMzMzMzMzMzMzMzMzMzNERERERERERERmZmZVVVVVVVVVVVVERERERERERERERERERERVVVVmZmZERERVVVVERERERERERERERERERERERERERERVVVVVVVVERERERERVVVVmZmZmZmZVVVVmZmZVVVVmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVERERVVVVVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZVVVVmZmZmZmZVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZVVVVVVVVmZmZVVVVmZmZmZmZ3d3dmZmZ3d3d3d3eIiIh3d3d3d3eIiIiIiIiIiIiIiIiIiIiZmZmZmZmIiIiZmZmIiIiIiIiZmZmZmZmqqqq7u7u7u7u7u7vMzMzMzMzd3d3d3d3d3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u3d3d3d3dzMzMzMzMqqqqqqqqmZmZmZmZqqqqqqqqqqqqqqqqqqqqqqqqqqqqu7u7qqqqqqqqmZmZmZmZqqqqmZmZmZmZmZmZqqqqqqqqqqqqqqqqqqqqqqqqmZmZmZmZmZmZmZmZd3d3iIiIiIiId3d3d3d3d3d3ZmZmVVVVREREREREMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREREREREREREREREREREREREREMzMzMzMzREREMzMzREREMzMzMzMzMzMzMzMzMzMzVVVVVVVVREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREREREREREREREREREVVVVVVVVVVVVREREVVVVREREREREVVVVREREVVVVREREVVVVVVVVVVVVZmZmZmZmVVVVZmZmZmZmd3d3d3d3ZmZmZmZmZmZmZmZmd3d3ZmZmZmZmVVVVZmZmZmZmd3d3ZmZmd3d3d3d3iIiIZmZmZmZmZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmd3d3d3d3ZmZmVVVVVVVVVVVVVVVVREREVVVVREREREREREREVVVVVVVVVVVVZmZmZmZmd3d3iIiIiIiImZmZiIiIiIiId3d3d3d3ZmZmZmZmVVVVZmZmZmZmZmZmiIiIiIiIiIiId3d3d3d3ZmZmZmZmZmZmZmZmVVVVZmZmZmZmd3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3iIiIiIiImZmZmZmZiIiImZmZd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiImZmZu7u7zMzMu7u7u7u7u7u7qqqqmZmZmZmZqqqqqqqqu7u7u7u7zMzM7u7uzMzMu7u7qqqqqqqqmZmZmZmZiIiIiIiIiIiImZmZmZmZqqqqmZmZiIiIiIiIqqqqmZmZqqqqqqqqmZmZmZmZmZmZmZmZqqqqqqqqqqqqqqqqu7u7qqqqqqqqqqqqqqqqmZmZqqqqu7u7u7u7u7u7qqqqqqqqqqqqqqqqmZmZmZmZmZmZmZmZmZmZiIiImZmZmZmZmZmZiIiIiIiImZmZmZmZqqqqmZmZmZmZmZmZmZmZiIiIiIiIiIiIiIiIiIiId3d3mZmZiIiId3d3d3d3iIiIiIiIiIiIqqqqqqqqqqqqmZmZmZmZmZmZiIiIiIiIiIiId3d3mZmZqqqqmZmZmZmZu7u7u7u7zMzMu7u7u7u7u7u7u7u7qqqqu7u7qqqqqqqqqqqqmZmZmZmZmZmZmZmZiIiIiIiIiIiId3d3d3d3ZmZmd3d3ZmZmZmZmVVVVZmZmVVVVZmZmVVVVVVVVZmZmVVVVVVVVREREREREVVVVREREVVVVREREMzMzMzMzREREMzMzREREREREMzMzREREMzMzREREMzMzMzMzMzMzMzMzMzMzIiIiIiIiIiIiIiIiIiIiMzMzIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiMzMzIiIiMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzMzMzREREMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREMzMzREREREREVVVVVVVVVVVVZmZmZmZmVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVVVVVREREREREREREREREREREVVVVVVVVVVVVVVVVZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3ZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3ZmZmd3d3d3d3d3d3ZmZmd3d3d3d3d3d3ZmZmZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3ZmZmd3d3d3d3iIiImZmZmZmZmZmZmZmZmZmZmZmZqqqqqqqqu7u7u7u7u7u7zMzMu7u7u7u7u7u7u7u7zMzM3d3d3d3d3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7szMzKqqqpmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmaqqqpmZmZmZmYiIiJmZmYiIiIiIiIiIiIiIiHd3d4iIiHd3d3d3d2ZmZmZmZlVVVVVVVVVVVWZmZlVVVVVVVWZmZlVVVVVVVURERFVVVURERERERDMzM0RERERERDMzMzMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERDMzMzMzM0RERERERERERERERERERERERERERERERDMzMzMzMzMzMzMzM0RERDMzM0RERERERERERERERERERERERERERERERERERERERERERERERERERDMzMzMzMzMzMzMzMyIiIjMzMzMzMzMzM2ZmZlVVVURERERERERERERERERERDMzMzMzM0RERERERERERERERFVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZlVVVVVVVXd3d2ZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d2ZmZmZmZlVVVWZmZmZmZmZmZnd3d3d3d3d3d3d3d4iIiHd3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d2ZmZnd3d3d3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVWZmZnd3d3d3d4iIiIiIiJmZmYiIiIiIiIiIiHd3d2ZmZmZmZmZmZmZmZmZmZnd3d4iIiIiIiJmZmYiIiIiIiHd3d1VVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d3d3d4iIiJmZmYiIiJmZmYiIiIiIiIiIiHd3d3d3d3d3d4iIiJmZmYiIiJmZmYiIiIiIiHd3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiKqqqqqqqru7u93d3e7u7u7u7t3d3e7u7t3d3czMzMzMzLu7u7u7u8zMzMzMzO7u7u7u7v///////93d3d3d3czMzKqqqqqqqpmZmZmZmaqqqqqqqpmZmaqqqqqqqqqqqpmZmZmZmZmZmZmZmaqqqqqqqpmZmZmZmaqqqru7u7u7u7u7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqru7u7u7u7u7u7u7u7u7u7u7u6qqqru7u6qqqpmZmZmZmZmZmZmZmZmZmaqqqqqqqpmZmZmZmZmZmaqqqpmZmaqqqqqqqpmZmYiIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiJmZmZmZmYiIiJmZmYiIiJmZmZmZmaqqqqqqqqqqqpmZmaqqqpmZmZmZmYiIiIiIiIiIiJmZmaqqqqqqqqqqqqqqqru7u8zMzLu7u8zMzLu7u6qqqqqqqqqqqqqqqqqqqpmZmZmZmZmZmZmZmYiIiIiIiHd3d3d3d3d3d2ZmZmZmZlVVVVVVVVVVVVVVVVVVVURERERERFVVVURERERERFVVVURERERERDMzM0RERERERDMzMzMzMzMzMzMzMzMzMzMzMzMzMyIiIiIiIiIiIiIiIiIiIiIiIiIiIjMzMyIiIiIiIiIiIiIiIiIiIjMzMzMzMyIiIjMzMyIiIiIiIjMzMzMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzMyIiIjMzM0RERERERERERDMzMzMzMzMzMzMzMzMzM0RERDMzM0RERERERFVVVVVVVURERFVVVWZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZlVVVVVVVWZmZmZmZnd3d2ZmZmZmZlVVVVVVVVVVVURERFVVVVVVVWZmZnd3d3d3d3d3d3d3d4iIiIiIiIiIiHd3d2ZmZmZmZmZmZlVVVVVVVWZmZmZmZnd3d2ZmZmZmZnd3d3d3d2ZmZnd3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d4iIiIiIiJmZmZmZmaqqqqqqqru7u7u7u8zMzMzMzMzMzN3d3d3d3d3d3e7u7u7u7u7u7u7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////u7u7d3d3MzMy7u7u7u7u7u7uqqqqZmZmIiIiIiIh3d3d3d3d3d3eIiIh3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3dmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3eIiIiIiIiIiIiIiIiZmZmIiIiZmZl3d3dERERVVVVEREREREQzMzNERERERERERERERERERERERERERERERERVVVVVVVVERERVVVVERERVVVVVVVVVVVVERERVVVVERERERERERERERERERERERERERERERERERERVVVVERERVVVVVVVVmZmZmZmZ3d3dVVVUzMzMzMzNEREREREQzMzMzMzMzMzNERERERER3d3d3d3dmZmZmZmZmZmZ3d3dmZmZVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3dmZmZ3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3dmZmZ3d3eIiIh3d3dmZmaIiIiIiIh3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3dmZmZ3d3d3d3eIiIiIiIh3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3dmZmZ3d3dmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZ3d3d3d3eIiIiIiIiZmZmIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3dmZmZ3d3d3d3eIiIiIiIiZmZmqqqqqqqqqqqqZmZmIiIh3d3dVVVVVVVVmZmZmZmZ3d3d3d3d3d3eZmZmIiIiZmZmZmZmZmZmZmZmZmZmIiIiIiIiIiIiIiIh3d3eIiIiIiIiZmZmZmZmZmZmqqqqIiIiIiIiIiIiIiIiIiIiZmZm7u7vMzMzd3d3u7u7////////////////////////////////u7u7u7u7d3d3d3d3u7u7////////////////////////////u7u7d3d3MzMzMzMzMzMzd3d3MzMzMzMy7u7u7u7u7u7u7u7uqqqqqqqqqqqqqqqqqqqqZmZmqqqqqqqq7u7u7u7u7u7uqqqqqqqqqqqqZmZmqqqqqqqqqqqq7u7u7u7uqqqq7u7u7u7uqqqqqqqqqqqqZmZmZmZmIiIiIiIiIiIiZmZmZmZmqqqqZmZmqqqqqqqqqqqqqqqqqqqqZmZmZmZmZmZmqqqqZmZmIiIiIiIiIiIiIiIiIiIiZmZmZmZmZmZmIiIiZmZmZmZmZmZmIiIiIiIiZmZmIiIiZmZmZmZmIiIiIiIiIiIiIiIiZmZmZmZmZmZmZmZmqqqqqqqqqqqq7u7u7u7u7u7uZmZmZmZmZmZmZmZmZmZmIiIiIiIiIiIiIiIiIiIiIiIh3d3dmZmZmZmZmZmZVVVVVVVVVVVVEREREREQzMzMzMzNEREQzMzNEREQzMzMzMzNEREQzMzMzMzMzMzMzMzMiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIzMzMiIiIiIiIzMzMzMzNEREREREREREREREREREREREREREREREQzMzNEREQzMzNEREREREQzMzMzMzMzMzMzMzMzMzMzMzMzMzMiIiIiIiIzMzMzMzMzMzMiIiIzMzMzMzNEREREREQzMzMzMzMzMzMzMzMzMzNERERERERVVVVVVVVmZmZ3d3d3d3dmZmZmZmZ3d3d3d3d3d3eIiIiIiIiIiIh3d3d3d3d3d3dmZmZ3d3d3d3d3d3eIiIh3d3d3d3dmZmZ3d3dmZmZmZmZmZmZmZmZ3d3d3d3d3d3dmZmZ3d3dmZmZ3d3d3d3dmZmZmZmZ3d3dmZmZ3d3dmZmZmZmZ3d3d3d3d3d3eIiIh3d3d3d3eIiIh3d3eIiIh3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3eIiIiZmZmZmZmZmZmZmZm7u7u7u7vMzMzd3d3d3d3d3d3u7u7u7u7u7u7////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3d3d3dzMzMu7u7u7u7qqqqmZmZqqqqqqqqqqqqmZmZmZmZmZmZqqqqqqqqqqqqu7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqqqqqqqqqu7u7u7u7u7u7u7u7u7u7u7u7qqqqmZmZiIiIZmZmREREVVVVREREREREREREREREREREREREREREREREVVVVREREVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVVVVVZmZmd3d3d3d3iIiImZmZmZmZqqqqu7u7qqqqZmZmREREMzMzZmZmZmZmREREMzMzREREVVVVZmZmd3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3iIiId3d3iIiId3d3iIiId3d3d3d3d3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3ZmZmd3d3ZmZmd3d3d3d3d3d3d3d3d3d3d3d3ZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3iIiImZmZmZmZmZmZmZmZmZmZiIiIiIiIiIiId3d3iIiIiIiIiIiIiIiIiIiImZmZqqqqqqqqu7u7u7u7u7u7qqqqqqqqqqqqiIiIiIiIZmZmd3d3d3d3d3d3iIiIiIiImZmZqqqqmZmZmZmZmZmZmZmZiIiImZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZqqqqqqqqqqqqmZmZmZmZiIiIiIiIqqqqu7u7zMzM7u7u7u7u////////////////////////////////////////////////7u7u////////////////////////////////////////////////7u7u////////7u7u7u7u7u7u7u7u7u7u7u7u3d3dzMzMzMzMu7u7u7u7u7u7u7u7u7u7zMzMu7u7u7u7qqqqu7u7qqqqqqqqu7u7u7u7qqqqu7u7qqqqu7u7qqqqqqqqqqqqmZmZqqqqmZmZiIiImZmZiIiImZmZmZmZmZmZmZmZqqqqqqqqu7u7qqqqu7u7qqqqqqqqmZmZmZmZiIiImZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZiIiImZmZmZmZmZmZqqqqqqqqu7u7qqqqqqqqmZmZmZmZiIiIiIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3ZmZmVVVVVVVVVVVVREREREREREREREREREREMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzMzMzMzMzMzMzIiIiMzMzIiIiMzMzMzMzMzMzREREREREREREREREREREREREMzMzREREVVVVZmZmZmZmZmZmZmZmd3d3ZmZmd3d3ZmZmVVVVVVVVREREREREREREREREREREMzMzMzMzREREMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzREREVVVVVVVVVVVVREREVVVVZmZmZmZmd3d3d3d3iIiIiIiIiIiId3d3iIiId3d3iIiImZmZiIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3iIiId3d3d3d3d3d3d3d3iIiId3d3iIiId3d3iIiId3d3d3d3d3d3d3d3iIiId3d3d3d3d3d3iIiIiIiId3d3iIiId3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZmZmZqqqqqqqqu7u7u7u7zMzM3d3dzMzM3d3d3d3d3d3d7u7u7u7u////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7t3d3d3d3czMzMzMzMzMzLu7u8zMzLu7u7u7u7u7u7u7u7u7u7u7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqoiIiHd3d2ZmZmZmZmZmZlVVVURERERERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVURERERERERERFVVVVVVVVVVVWZmZlVVVWZmZnd3d3d3d3d3d4iIiGZmZnd3d4iIiJmZmaqqqru7u7u7u8zMzMzMzMzMzMzMzN3d3czMzIiIiERERERERGZmZmZmZkRERERERERERGZmZnd3d3d3d2ZmZnd3d2ZmZnd3d3d3d2ZmZmZmZmZmZnd3d3d3d4iIiHd3d3d3d3d3d2ZmZoiIiIiIiIiIiHd3d4iIiIiIiJmZmYiIiIiIiHd3d3d3d2ZmZnd3d3d3d4iIiHd3d3d3d3d3d3d3d2ZmZnd3d2ZmZmZmZnd3d2ZmZmZmZnd3d3d3d4iIiHd3d3d3d3d3d3d3d4iIiHd3d3d3d3d3d2ZmZnd3d2ZmZmZmZmZmZnd3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiIiIiJmZmZmZmZmZmZmZmaqqqqqqqpmZmaqqqoiIiJmZmYiIiIiIiHd3d4iIiIiIiJmZmaqqqru7u7u7u8zMzLu7u8zMzLu7u7u7u6qqqqqqqpmZmZmZmYiIiIiIiHd3d3d3d4iIiJmZmZmZmaqqqqqqqpmZmYiIiIiIiIiIiIiIiIiIiJmZmZmZmZmZmZmZmaqqqpmZmZmZmaqqqpmZmaqqqru7u6qqqpmZmYiIiJmZmaqqqszMzO7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////+7u7t3d3e7u7t3d3czMzLu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqqqqqpmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiJmZmaqqqqqqqqqqqru7u6qqqru7u7u7u6qqqqqqqoiIiIiIiJmZmYiIiIiIiHd3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d3d3d4iIiIiIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiKqqqqqqqqqqqru7u6qqqru7u6qqqpmZmZmZmXd3d3d3d3d3d2ZmZlVVVWZmZlVVVVVVVVVVVVVVVVVVVURERERERDMzM0RERDMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzM0RERERERDMzM0RERERERERERERERERERERERFVVVVVVVWZmZnd3d2ZmZmZmZmZmZlVVVVVVVVVVVWZmZmZmZnd3d2ZmZmZmZnd3d3d3d3d3d3d3d2ZmZlVVVVVVVURERERERERERERERERERERERDMzM0RERDMzMzMzM0RERERERERERDMzM0RERERERERERERERDMzM0RERERERGZmZmZmZmZmZmZmZmZmZmZmZnd3d4iIiHd3d4iIiIiIiJmZmYiIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d4iIiIiIiHd3d3d3d3d3d3d3d4iIiIiIiIiIiIiIiIiIiJmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiJmZmYiIiIiIiIiIiHd3d4iIiIiIiIiIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiKqqqqqqqqqqqqqqqru7u8zMzMzMzN3d3d3d3e7u7u7u7u7u7v///////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3d3d3d3d3d3d3d3d27u7u7u7u7u7uqqqqqqqqqqqqZmZmZmZmZmZmZmZmZmZmqqqqqqqqqqqqqqqqZmZl3d3dmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3eIiIiIiIiZmZmZmZmIiIh3d3d3d3dmZmZ3d3eIiIiZmZmZmZmqqqqqqqq7u7vMzMzMzMzMzMzMzMy7u7vMzMzd3d3d3d3d3d3d3d3MzMzd3d3d3d3d3d3d3d3d3d2qqqpmZmZERER3d3eIiIhVVVUzMzNERERmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZ3d3eIiIiZmZmZmZmIiIiZmZmIiIiZmZmIiIiIiIiIiIh3d3d3d3dmZmZ3d3d3d3eIiIh3d3d3d3dmZmZ3d3dmZmZmZmZ3d3d3d3dmZmZ3d3d3d3eIiIiIiIiIiIh3d3d3d3d3d3eIiIh3d3dmZmZ3d3dmZmZ3d3dmZmZ3d3d3d3eIiIiIiIiZmZmZmZmZmZmqqqqqqqqqqqq7u7uqqqqqqqqqqqqqqqq7u7uqqqq7u7uqqqqqqqqZmZmZmZmIiIiIiIiZmZmqqqqqqqq7u7vMzMy7u7vMzMy7u7u7u7u7u7uqqqqqqqqZmZmZmZmqqqqZmZmIiIiZmZmIiIiIiIiZmZmqqqqZmZmZmZmIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZmZmZmZmZmqqqq7u7uqqqqqqqq7u7u7u7uqqqqZmZmqqqqqqqq7u7vd3d3////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////u7u7u7u7d3d3MzMy7u7u7u7u7u7u7u7u7u7vMzMy7u7u7u7uqqqq7u7uqqqqZmZmZmZmZmZmqqqqqqqqqqqqqqqqZmZmZmZmZmZmqqqq7u7u7u7u7u7u7u7u7u7uqqqqqqqqqqqqZmZmIiIiIiIiIiIiIiIh3d3eIiIh3d3d3d3eIiIh3d3d3d3d3d3d3d3eIiIh3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZl3d3eIiIiIiIiZmZmqqqqqqqqqqqqqqqqqqqqqqqqqqqqIiIiIiIh3d3dmZmZVVVVVVVVVVVVERERERERVVVVEREQzMzNERERVVVVVVVVERERERERERERERERVVVVERERVVVVVVVVVVVVmZmZ3d3dmZmZmZmZmZmZmZmZmZmZVVVVVVVVVVVVmZmZmZmZ3d3eIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERVVVVERERVVVVVVVVVVVVVVVVERERVVVVmZmZVVVVVVVVVVVVmZmZVVVVVVVVVVVVERERmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIh3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiZmZmZmZmZmZmIiIiZmZmIiIiZmZmIiIiIiIiZmZmZmZmIiIiZmZmIiIiIiIiZmZmZmZmIiIiIiIiIiIiZmZmZmZmqqqqZmZmZmZmZmZmZmZmIiIiZmZmqqqqqqqq7u7u7u7u7u7vMzMzd3d3d3d3u7u7u7u7////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7///////////////////8A//8AAP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7d3d3d3d3d3d3d3d27u7u7u7u7u7u7u7vMzMzd3d3d3d3d3d3d3d3MzMy7u7uqqqqZmZmqqqqqqqq7u7uqqqq7u7u7u7u7u7vMzMzMzMzd3d3d3d3u7u7u7u7u7u7u7u7u7u7d3d3d3d3MzMzd3d3d3d3u7u7u7u7u7u7////u7u7////u7u7////u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3d3d3d3d3u7u67u7uIiIhmZmZmZmZ3d3dVVVVERERmZmZ3d3eIiIh3d3dmZmZ3d3dmZmZ3d3d3d3d3d3d3d3dmZmZmZmZVVVVVVVVmZmZ3d3d3d3eIiIiIiIiIiIiIiIiIiIiZmZmIiIiIiIiIiIh3d3eIiIh3d3eIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3d3d3eZmZmIiIiIiIh3d3d3d3d3d3d3d3eIiIiIiIiIiIiZmZmZmZmZmZmqqqqZmZmqqqqqqqqqqqqZmZmqqqqqqqq7u7u7u7u7u7u7u7u7u7vMzMy7u7u7u7vMzMy7u7u7u7u7u7uqqqqqqqq7u7u7u7vMzMzd3d3MzMzMzMy7u7u7u7u7u7uqqqqqqqqqqqqZmZmqqqqqqqqqqqqZmZmZmZmqqqqZmZmqqqqZmZmIiIh3d3d3d3d3d3eIiIiIiIiZmZmZmZmqqqqqqqqqqqqqqqq7u7uqqqq7u7uqqqq7u7uqqqqqqqqqqqqqqqrMzMzd3d3u7u7////////////////////////////////////////u7u7////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////u7u7d3d3MzMzMzMy7u7vMzMy7u7u7u7u7u7u7u7uqqqqqqqqqqqqqqqqqqqqZmZmqqqqZmZmZmZmqqqqZmZmqqqqqqqqqqqq7u7u7u7u7u7uqqqqqqqqZmZmZmZmIiIiIiIiIiIiIiIh3d3eIiIiIiIiIiIiIiIh3d3d3d3eIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3eIiIh3d3d3d3d3d3eIiIh3d3eIiIiIiIiIiIh3d3d3d3dmZmZmZmZVVVVEREREREREREQzMzMzMzMiIiIzMzMzMzNEREQzMzNERERERERmZmZmZmZ3d3dmZmZVVVVmZmZmZmZ3d3d3d3eIiIiIiIiZmZmqqqqZmZmZmZmIiIh3d3d3d3d3d3d3d3eIiIh3d3eIiIiZmZmIiIiZmZmIiIiIiIh3d3eIiIiIiIh3d3eIiIh3d3d3d3d3d3d3d3dmZmZVVVVVVVVVVVVmZmZVVVVERERVVVVERERmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3dmZmZ3d3d3d3d3d3d3d3dmZmZ3d3d3d3dmZmZ3d3d3d3d3d3d3d3eIiIiIiIh3d3eIiIiIiIiIiIiIiIiIiIiZmZmIiIiIiIiIiIiIiIiZmZmZmZmIiIiZmZmIiIiZmZmZmZmIiIh3d3d3d3d3d3eIiIiZmZmIiIiIiIiZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmqqqqqqqqZmZmZmZmZmZmZmZmZmZmZmZmZmZmqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqq7u7vMzMzMzMzd3d3d3d3u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u////////7u7u////////////7u7u////7u7u////7u7u////////7u7u////////////////////////////////////////////////////////////////////////7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3dqqqqZmZmZmZmZmZmREREVVVVd3d3d3d3d3d3ZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmVVVVVVVVREREVVVVZmZmd3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiId3d3d3d3d3d3iIiId3d3iIiId3d3d3d3d3d3ZmZmd3d3d3d3iIiImZmZiIiIqqqqqqqqqqqqqqqqu7u7qqqqu7u7qqqqqqqqqqqqqqqqmZmZmZmZqqqqqqqqu7u7u7u7u7u7u7u7u7u7u7u7zMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7zMzMzMzMzMzMzMzMu7u7u7u7u7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqqqqqu7u7qqqqqqqqqqqqqqqqqqqqmZmZiIiId3d3d3d3iIiImZmZqqqqqqqqu7u7u7u7zMzMu7u7zMzMu7u7zMzMu7u7qqqqu7u7u7u7u7u7qqqqzMzM3d3d7u7u////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////3d3d3d3dzMzMzMzMzMzMu7u7u7u7u7u7u7u7u7u7qqqqqqqqmZmZqqqqmZmZqqqqqqqqmZmZqqqqmZmZqqqqqqqqmZmZqqqqmZmZqqqqmZmZmZmZiIiIiIiIiIiId3d3iIiId3d3iIiIiIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3ZmZmVVVVZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREVVVVREREREREREREMzMzREREREREREREMzMzMzMzMzMzMzMzIiIiMzMzMzMzMzMzMzMzREREREREVVVVZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiImZmZiIiIiIiId3d3d3d3d3d3iIiId3d3iIiIiIiIiIiIiIiId3d3iIiIiIiIiIiId3d3d3d3d3d3iIiId3d3iIiIiIiId3d3d3d3d3d3ZmZmd3d3ZmZmZmZmd3d3ZmZmZmZmZmZmd3d3d3d3d3d3d3d3iIiIiIiIiIiId3d3iIiId3d3d3d3iIiIiIiId3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZmZmZiIiImZmZiIiImZmZiIiIiIiImZmZmZmZmZmZmZmZmZmZiIiIiIiId3d3iIiIiIiIiIiIiIiImZmZmZmZmZmZmZmZmZmZmZmZmZmZiIiImZmZiIiId3d3iIiIiIiImZmZmZmZmZmZmZmZmZmZmZmZmZmZqqqqu7u7zMzMu7u7u7u7u7u7u7u7u7u7zMzM3d3d3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7u7u7t3d3d3d3d3d3czMzN3d3czMzMzMzMzMzMzMzMzMzMzMzMzMzN3d3czMzLu7u3d3d2ZmZlVVVVVVVWZmZmZmZlVVVVVVVWZmZlVVVVVVVVVVVWZmZmZmZnd3d3d3d2ZmZmZmZnd3d3d3d4iIiIiIiIiIiJmZmZmZmZmZmYiIiIiIiHd3d3d3d3d3d2ZmZnd3d2ZmZnd3d3d3d4iIiIiIiHd3d3d3d3d3d4iIiHd3d4iIiIiIiIiIiHd3d4iIiIiIiIiIiIiIiJmZmZmZmZmZmaqqqru7u7u7u7u7u7u7u6qqqqqqqqqqqpmZmZmZmZmZmaqqqqqqqqqqqru7u7u7u8zMzMzMzMzMzLu7u7u7u7u7u8zMzLu7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqqqqqru7u6qqqqqqqru7u6qqqru7u6qqqru7u7u7u7u7u6qqqqqqqqqqqqqqqpmZmZmZmZmZmYiIiJmZmaqqqru7u7u7u8zMzN3d3d3d3czMzMzMzMzMzMzMzKqqqqqqqqqqqru7u93d3czMzO7u7u7u7v///////////////////////////////////////+7u7v///////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////+7u7v///////////////////+7u7v///////////////////////+7u7v///////////+7u7t3d3czMzMzMzMzMzLu7u7u7u7u7u7u7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqpmZmaqqqpmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiIiIiHd3d3d3d3d3d2ZmZnd3d2ZmZnd3d2ZmZmZmZmZmZlVVVVVVVVVVVURERERERERERERERERERFVVVURERERERFVVVURERFVVVVVVVVVVVVVVVURERDMzM0RERERERERERERERERERFVVVVVVVVVVVURERERERDMzM0RERDMzM0RERDMzM0RERFVVVVVVVXd3d3d3d4iIiHd3d4iIiIiIiHd3d3d3d3d3d2ZmZnd3d2ZmZmZmZnd3d4iIiGZmZnd3d2ZmZmZmZmZmZnd3d2ZmZnd3d4iIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiHd3d3d3d3d3d3d3d3d3d3d3d4iIiHd3d4iIiHd3d4iIiHd3d4iIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d4iIiIiIiIiIiIiIiIiIiHd3d4iIiIiIiIiIiJmZmZmZmZmZmYiIiJmZmaqqqqqqqpmZmaqqqqqqqqqqqpmZmZmZmZmZmZmZmZmZmYiIiJmZmYiIiIiIiJmZmYiIiJmZmYiIiJmZmYiIiIiIiIiIiJmZmYiIiIiIiIiIiHd3d3d3d3d3d4iIiIiIiJmZmZmZmZmZmZmZmZmZmaqqqqqqqqqqqru7u7u7u7u7u7u7u8zMzN3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3d3d3MzMzMzMzMzMy7u7u7u7uqqqqqqqqqqqq7u7u7u7u7u7u7u7uIiIhmZmZVVVVmZmZmZmZVVVVVVVVVVVVmZmZmZmZmZmZ3d3eIiIiIiIiZmZmZmZmqqqqZmZmqqqqqqqq7u7u7u7uqqqqZmZmZmZmIiIiIiIh3d3dmZmZmZmZmZmZmZmZ3d3dmZmZmZmZ3d3d3d3d3d3d3d3eZmZmIiIiZmZmZmZmZmZmZmZmqqqq7u7uqqqq7u7u7u7vMzMy7u7u7u7uqqqqqqqq7u7uqqqqqqqqqqqqqqqqqqqqZmZmqqqqqqqq7u7u7u7u7u7vMzMy7u7vMzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7uqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqZmZmqqqqqqqqqqqq7u7u7u7u7u7u7u7uqqqq7u7u7u7u7u7vMzMzMzMyqqqqqqqqqqqqqqqq7u7u7u7vMzMzMzMzMzMzMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d27u7u7u7u7u7uqqqq7u7vMzMzu7u7u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////u7u7u7u7u7u7d3d3u7u7d3d3MzMzd3d3d3d3d3d3d3d3d3d3d3d3d3d3MzMy7u7u7u7uZmZmZmZmIiIiIiIiIiIiZmZmIiIh3d3dmZmZ3d3dmZmZmZmZmZmZVVVVVVVVmZmZ3d3dmZmZERERVVVVERERERERVVVVVVVVVVVVVVVVERERmZmZVVVVmZmZmZmZVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmaIiIiIiIiIiIhmZmZVVVVmZmZmZmZmZmZ3d3dmZmZ3d3eIiIiZmZmZmZmZmZmqqqqZmZmqqqqZmZmIiIh3d3d3d3d3d3d3d3dmZmZ3d3eIiIh3d3dmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3eIiIh3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIh3d3d3d3d3d3eIiIh3d3eIiIiIiIh3d3eIiIh3d3eIiIiIiIiIiIiIiIiZmZmIiIiIiIiIiIiIiIiIiIiZmZmZmZmqqqqZmZmZmZmZmZmZmZmqqqqZmZmqqqqZmZmqqqqqqqqqqqqqqqqqqqqZmZmqqqqZmZmqqqqqqqq7u7uqqqqqqqqZmZmZmZmqqqqqqqqqqqqZmZmZmZmZmZmqqqqZmZmZmZmZmZmIiIiIiIiIiIh3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3eIiIh3d3eIiIiIiIiIiIiIiIiIiIiqqqqqqqq7u7uqqqq7u7u7u7vMzMzd3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////7u7u7u7u7u7u3d3d3d3dzMzMzMzMu7u7u7u7u7u7u7u7qqqqu7u7qqqqiIiId3d3d3d3ZmZmZmZmZmZmiIiImZmZmZmZmZmZmZmZmZmZqqqqu7u7qqqqu7u7u7u7u7u7u7u7u7u7qqqqmZmZmZmZiIiImZmZd3d3d3d3ZmZmd3d3d3d3d3d3ZmZmd3d3d3d3d3d3d3d3iIiIqqqqu7u7zMzMzMzMzMzMzMzMzMzM3d3dzMzM3d3d3d3dzMzMzMzMzMzMu7u7u7u7zMzMu7u7zMzMu7u7u7u7u7u7qqqqu7u7u7u7u7u7u7u7zMzMzMzMu7u7u7u7u7u7u7u7u7u7u7u7u7u7qqqqqqqqqqqqmZmZmZmZiIiImZmZiIiIqqqqqqqqu7u7qqqqu7u7u7u7u7u7u7u7qqqqqqqqqqqqqqqqu7u7u7u7u7u7u7u7zMzMzMzMu7u7u7u7u7u7zMzM3d3d3d3d3d3d7u7u3d3d7u7u3d3d3d3dzMzMzMzMzMzMu7u7zMzMu7u7zMzMzMzM3d3d////////////////////////////////////////////////7u7u////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////7u7u////////////////////////////////////////7u7u////////////////7u7u3d3dzMzMu7u7qqqqqqqqiIiIiIiIiIiIiIiId3d3ZmZmZmZmd3d3d3d3mZmZd3d3ZmZmVVVVVVVVZmZmVVVVZmZmZmZmd3d3ZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3iIiId3d3ZmZmZmZmd3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREREREREREVVVVREREVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVZmZmZmZmd3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmd3d3ZmZmZmZmd3d3d3d3d3d3d3d3d3d3iIiIiIiImZmZmZmZmZmZqqqqqqqqu7u7qqqqu7u7qqqqqqqqqqqqqqqqqqqqqqqqqqqqmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZiIiImZmZiIiIiIiIiIiIiIiId3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3iIiId3d3mZmZmZmZqqqqqqqqu7u7qqqqu7u7zMzMzMzM3d3d////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7t3d3e7u7t3d3d3d3d3d3czMzLu7u6qqqpmZmaqqqqqqqqqqqru7u6qqqru7u8zMzMzMzMzMzLu7u6qqqqqqqqqqqru7u6qqqqqqqpmZmYiIiIiIiIiIiJmZmYiIiIiIiIiIiJmZmYiIiJmZmYiIiJmZmaqqqqqqqru7u8zMzN3d3d3d3e7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3czMzMzMzMzMzMzMzMzMzN3d3czMzN3d3d3d3czMzLu7u7u7u8zMzLu7u7u7u7u7u7u7u7u7u6qqqru7u6qqqru7u6qqqqqqqqqqqpmZmaqqqpmZmZmZmZmZmZmZmaqqqru7u8zMzN3d3d3d3d3d3czMzLu7u7u7u5mZmYiIiJmZmZmZmaqqqru7u7u7u7u7u8zMzMzMzMzMzMzMzMzMzMzMzN3d3d3d3e7u7u7u7u7u7u7u7u7u7t3d3d3d3czMzMzMzMzMzMzMzMzMzMzMzO7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////+7u7v///////////////////////////////93d3czMzLu7u6qqqpmZmZmZmZmZmZmZmZmZmYiIiHd3d3d3d3d3d3d3d4iIiHd3d3d3d3d3d2ZmZmZmZnd3d3d3d3d3d3d3d2ZmZmZmZnd3d2ZmZlVVVVVVVVVVVURERFVVVURERERERFVVVVVVVURERERERERERFVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVURERFVVVVVVVWZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZlVVVVVVVURERFVVVURERFVVVURERERERERERERERERERERERFVVVURERERERFVVVVVVVVVVVVVVVWZmZnd3d2ZmZnd3d3d3d3d3d2ZmZmZmZmZmZmZmZlVVVURERERERFVVVVVVVVVVVWZmZmZmZnd3d4iIiIiIiIiIiJmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmYiIiIiIiHd3d3d3d3d3d3d3d3d3d2ZmZnd3d2ZmZmZmZmZmZlVVVWZmZlVVVVVVVWZmZlVVVVVVVVVVVURERFVVVURERERERERERERERERERFVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d4iIiIiIiJmZmZmZmaqqqru7u7u7u7u7u7u7u7u7u8zMzN3d3d3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3u7u7u7u7////u7u7d3d3MzMzMzMzd3d3d3d3MzMzMzMy7u7uqqqq7u7uqqqqqqqq7u7uqqqq7u7u7u7vMzMzMzMzd3d3d3d3u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3d3d3MzMzd3d3d3d3MzMzd3d3d3d3d3d27u7u7u7u7u7u7u7u7u7u7u7u7u7uqqqqqqqqqqqqZmZmqqqqqqqqZmZmZmZmZmZmZmZmqqqqqqqq7u7vMzMzMzMzd3d3u7u7u7u7u7u7u7u7u7u7d3d27u7uqqqqIiIiIiIiZmZmZmZmqqqq7u7u7u7vMzMzMzMzd3d3d3d3d3d3d3d3d3d3d3d3u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3MzMzMzMzMzMzd3d3u7u7u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////u7u7u7u7////////////////////////////////////////////////////////////////////////////////u7u7////u7u7MzMyqqqqZmZmqqqqZmZmIiIiIiIiIiIh3d3eIiIiIiIhmZmZmZmZ3d3dmZmZVVVVmZmZVVVVmZmZmZmZmZmZmZmZ3d3dmZmZmZmZmZmZmZmZVVVVVVVVERERVVVVERERERERERERERERERERVVVVEREREREREREREREREREREREREREQzMzNERERERERERERERERERERERERERERERERERERERERERERERERERERERERVVVVERERVVVVERERERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVERERERERVVVVVVVVVVVVERERVVVVVVVVmZmZmZmZmZmZ3d3d3d3d3d3eIiIiIiIiIiIiIiIh3d3dmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3eIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3dmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVVVVVERERERERERERERERERERERERVVVVEREREREQzMzNERERERERERERVVVVERERVVVVmZmZmZmZ3d3d3d3d3d3eIiIiIiIiZmZmZmZmqqqq7u7u7u7u7u7u7u7vMzMzMzMzMzMzd3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u////7u7u////7u7u////7u7u////7u7u////7u7u3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMu7u7u7u7zMzMu7u7u7u7qqqqiIiImZmZqqqqqqqqqqqqqqqqmZmZqqqqmZmZmZmZmZmZmZmZmZmZqqqqqqqqu7u7zMzM3d3d7u7u7u7u////////////////////7u7u3d3dzMzMu7u7qqqqiIiImZmZmZmZqqqqu7u7qqqqzMzM3d3d7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d7u7u3d3d3d3d3d3dzMzM7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u////////////////////////7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3d3d3d3d3dzMzMzMzMu7u7qqqqmZmZd3d3d3d3ZmZmZmZmVVVVZmZmVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmVVVVVVVVZmZmd3d3ZmZmd3d3ZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVREREVVVVVVVVREREREREREREREREREREMzMzREREVVVVREREREREREREREREVVVVREREREREREREVVVVZmZmVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVZmZmVVVVVVVVVVVVZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVREREREREREREMzMzREREREREREREREREREREREREREREREREREREREREREREREREVVVVVVVVZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiIiIiImZmZqqqqu7u7u7u7u7u7zMzMu7u7zMzM3d3d3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3czMzMzMzMzMzLu7u7u7u7u7u6qqqqqqqqqqqqqqqqqqqqqqqoiIiGZmZoiIiJmZmaqqqpmZmaqqqqqqqqqqqqqqqqqqqru7u8zMzMzMzO7u7u7u7u7u7v///////////////////////////////+7u7u7u7t3d3czMzMzMzLu7u5mZmZmZmaqqqru7u7u7u8zMzO7u7u7u7u7u7v///+7u7u7u7u7u7u7u7v///+7u7u7u7t3d3e7u7u7u7u7u7u7u7u7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7v///////////////////////+7u7u7u7t3d3czMzMzMzMzMzMzMzMzMzLu7u8zMzLu7u7u7u6qqqoiIiIiIiHd3d2ZmZlVVVVVVVVVVVVVVVURERFVVVVVVVVVVVURERERERERERGZmZmZmZlVVVWZmZmZmZnd3d4iIiHd3d2ZmZmZmZnd3d4iIiHd3d3d3d3d3d3d3d2ZmZlVVVWZmZmZmZlVVVVVVVURERERERFVVVURERGZmZnd3d2ZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZnd3d2ZmZmZmZnd3d2ZmZmZmZmZmZmZmZnd3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d2ZmZmZmZmZmZmZmZmZmZmZmZmZmZnd3d2ZmZnd3d3d3d3d3d3d3d3d3d4iIiHd3d3d3d3d3d3d3d4iIiJmZmZmZmZmZmYiIiHd3d3d3d2ZmZlVVVVVVVVVVVWZmZlVVVURERERERFVVVVVVVVVVVWZmZmZmZmZmZmZmZlVVVVVVVWZmZlVVVVVVVVVVVVVVVVVVVURERFVVVVVVVVVVVVVVVURERFVVVURERFVVVURERERERERERERERERERERERERERERERERERERERERERERERFVVVURERERERFVVVURERFVVVVVVVWZmZmZmZnd3d3d3d3d3d3d3d4iIiHd3d4iIiJmZmaqqqqqqqru7u7u7u8zMzMzMzLu7u8zMzN3d3d3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////u7u7////u7u7////u7u7u7u7u7u7u7u7d3d3d3d3MzMy7u7u7u7vMzMy7u7u7u7u7u7u7u7u7u7u7u7uqqqqqqqq7u7uZmZmIiIh3d3eZmZmqqqq7u7u7u7vMzMzMzMzu7u7u7u7u7u7u7u7////////////////////////////////////////u7u7u7u7u7u7u7u7d3d3d3d3d3d3MzMyqqqqZmZmqqqqqqqrMzMzd3d3u7u7////u7u7u7u7////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7u7u7u7u7////////////////u7u7u7u7u7u7d3d3d3d3u7u7d3d3d3d3u7u7d3d3MzMzMzMy7u7uZmZmZmZmIiIiIiIiIiIhmZmZVVVVVVVVVVVVVVVVVVVVVVVVVVVVERERERERVVVVmZmZVVVVmZmZ3d3eIiIiIiIiIiIiIiIiIiIiIiIiIiIh3d3eIiIiIiIiIiIh3d3d3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZ3d3eIiIiIiIiIiIh3d3dmZmZ3d3d3d3d3d3eIiIiIiIiIiIiIiIiIiIh3d3d3d3d3d3eIiIh3d3dmZmZ3d3dmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3eIiIiIiIiIiIh3d3eIiIiZmZmZmZmZmZmZmZmZmZmqqqq7u7uqqqqZmZmqqqqqqqqZmZmIiIiZmZmqqqqqqqqqqqqIiIhmZmZERERERERERERVVVVmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZVVVVVVVVmZmZVVVVERERVVVVERERVVVVERERVVVVERERVVVVVVVVVVVVVVVVEREREREREREREREREREREREREREREREQzMzNEREQzMzNERERERERERERVVVVVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIiZmZm7u7u7u7vMzMy7u7vMzMzMzMzMzMzMzMzd3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////7u7u////////////////////////////////////////////////////////////////////////////7u7u7u7u////7u7u3d3d3d3d7u7u7u7u7u7u7u7u3d3d7u7u7u7u7u7u7u7u7u7u3d3dzMzMzMzM3d3d7u7u////7u7u////////////////////////////////////////////////////////////7u7u7u7u7u7u3d3d7u7u7u7u7u7u3d3d3d3du7u7qqqqmZmZqqqqu7u7zMzM7u7u7u7u////7u7u7u7u////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u7u7u7u7u3d3du7u7qqqqiIiImZmZmZmZqqqqmZmZiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiImZmZmZmZqqqqqqqqqqqqmZmZmZmZmZmZqqqqqqqqmZmZmZmZmZmZmZmZiIiId3d3iIiId3d3iIiId3d3iIiImZmZu7u7qqqqqqqqiIiIiIiIiIiId3d3iIiIiIiIiIiImZmZmZmZmZmZiIiIiIiIiIiIiIiIiIiIZmZmZmZmVVVVVVVVVVVVZmZmZmZmd3d3ZmZmVVVVZmZmd3d3mZmZqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqu7u7u7u7u7u7qqqqqqqqqqqqmZmZiIiIiIiIqqqqu7u7u7u7mZmZd3d3ZmZmZmZmZmZmZmZmZmZmd3d3ZmZmZmZmVVVVVVVVREREREREREREREREREREREREVVVVREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVREREVVVVREREREREREREVVVVREREREREREREREREREREREREREREVVVVVVVVZmZmZmZmd3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiImZmZmZmZqqqqqqqqu7u7zMzMzMzMzMzMzMzMzMzM3d3d3d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7u7u7u7u7u7u7u7u7t3d3czMzJmZmYiIiKqqqszMzO7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////+7u7t3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////93d3czMzMzMzMzMzMzMzMzMzLu7u6qqqqqqqqqqqpmZmaqqqpmZmaqqqpmZmaqqqqqqqqqqqqqqqqqqqpmZmbu7u8zMzMzMzKqqqpmZmYiIiIiIiIiIiHd3d3d3d3d3d4iIiIiIiIiIiLu7u93d3czMzLu7u6qqqpmZmZmZmZmZmZmZmZmZmYiIiJmZmZmZmZmZmaqqqqqqqqqqqpmZmYiIiIiIiGZmZnd3d2ZmZlVVVWZmZmZmZnd3d3d3d1VVVVVVVVVVVXd3d5mZmbu7u8zMzLu7u8zMzMzMzKqqqoiIiKqqqru7u8zMzMzMzKqqqqqqqqqqqpmZmZmZmbu7u6qqqru7u7u7u6qqqoiIiHd3d2ZmZmZmZmZmZlVVVURERERERERERERERERERERERERERFVVVVVVVVVVVVVVVURERFVVVWZmZlVVVVVVVVVVVURERFVVVURERFVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVURERERERERERERERFVVVWZmZmZmZnd3d3d3d4iIiHd3d4iIiHd3d4iIiHd3d3d3d4iIiIiIiIiIiJmZmaqqqru7u7u7u7u7u8zMzMzMzMzMzMzMzMzMzN3d3d3d3e7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7d3d27u7uZmZm7u7vu7u7////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7d3d3d3d3u7u7////////////////////////////////////////////////////////////////////u7u7////d3d3d3d3d3d3d3d3MzMzMzMzMzMyqqqqqqqqZmZmqqqqZmZmZmZmqqqqqqqqqqqqZmZmqqqqZmZmZmZm7u7vMzMy7u7u7u7uZmZmIiIiIiIh3d3d3d3eIiIiIiIiZmZmZmZmZmZnMzMzd3d3MzMzMzMy7u7u7u7u7u7u7u7uqqqqqqqqqqqqZmZmqqqq7u7uqqqqqqqqqqqqqqqqZmZmIiIiIiIiIiIhmZmZmZmZ3d3d3d3eIiIh3d3dVVVVVVVVmZmZ3d3eqqqrd3d3d3d3MzMzMzMzMzMyIiIhmZmZ3d3e7u7vMzMzMzMy7u7uqqqqqqqqqqqq7u7u7u7u7u7vMzMy7u7uqqqp3d3dmZmZVVVVVVVVVVVVVVVVERERERERERERERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZVVVVVVVVVVVVVVVVmZmZmZmZ3d3d3d3eIiIh3d3eIiIh3d3eIiIh3d3d3d3eIiIiIiIiIiIiZmZmqqqq7u7u7u7u7u7vMzMzMzMzd3d3MzMzMzMzMzMzd3d3d3d3u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u3d3d3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u3d3dzMzM3d3d////////////////////////////////////////////////////////////////////////////7u7u7u7u3d3d7u7u3d3d7u7uzMzMu7u7u7u7qqqqqqqqqqqqqqqqmZmZmZmZqqqqmZmZmZmZmZmZqqqqzMzMu7u7qqqqmZmZmZmZiIiIiIiIiIiIiIiIiIiImZmZqqqqu7u73d3d3d3dzMzMzMzMu7u7u7u7u7u7u7u7qqqqu7u7u7u7zMzMzMzMu7u7zMzMu7u7u7u7qqqqqqqqqqqqmZmZiIiId3d3iIiIiIiIiIiIiIiId3d3ZmZmZmZmd3d3mZmZzMzM3d3d3d3dzMzMu7u7iIiIZmZmZmZmZmZmiIiI3d3d3d3dzMzMu7u7u7u7u7u7zMzMu7u7u7u7zMzM3d3dqqqqd3d3VVVVREREREREVVVVREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVZmZmZmZmd3d3iIiId3d3iIiIiIiIiIiIiIiId3d3iIiId3d3iIiImZmZmZmZqqqqu7u7u7u7zMzMzMzMzMzMzMzMzMzM3d3dzMzMzMzM7u7u7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7t3d3czMzN3d3e7u7v///////////////////////////////////////////////////////////////////////////+7u7v///////////+7u7t3d3czMzLu7u7u7u7u7u6qqqqqqqqqqqqqqqpmZmZmZmZmZmaqqqru7u7u7u7u7u6qqqqqqqqqqqpmZmZmZmaqqqpmZmaqqqru7u8zMzN3d3czMzMzMzLu7u7u7u7u7u7u7u6qqqru7u8zMzN3d3d3d3czMzMzMzMzMzMzMzLu7u8zMzLu7u6qqqqqqqpmZmZmZmYiIiJmZmYiIiIiIiHd3d3d3d2ZmZnd3d7u7u93d3czMzMzMzLu7u5mZmXd3d3d3d3d3d2ZmZnd3d6qqqszMzMzMzMzMzMzMzMzMzLu7u6qqqru7u8zMzMzMzKqqqmZmZkRERERERFVVVURERFVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVWZmZmZmZmZmZnd3d3d3d4iIiHd3d4iIiHd3d4iIiHd3d3d3d3d3d3d3d4iIiJmZmaqqqru7u8zMzMzMzMzMzN3d3d3d3d3d3czMzN3d3d3d3d3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////u7u7u7u7MzMzd3d3u7u7u7u7////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3d3d3MzMzMzMy7u7uqqqq7u7uqqqqqqqqqqqq7u7vMzMy7u7vMzMyqqqqqqqq7u7u7u7uZmZmZmZm7u7u7u7u7u7vMzMzMzMy7u7u7u7u7u7vMzMy7u7u7u7uqqqqqqqrMzMzMzMzMzMzd3d3d3d3MzMzMzMzMzMy7u7u7u7u7u7uqqqqZmZmZmZmIiIiIiIiIiIiIiIh3d3eIiIiIiIiZmZm7u7vMzMy7u7u7u7uZmZmIiIh3d3d3d3d3d3dmZmZ3d3d3d3eqqqq7u7vMzMzMzMy7u7uqqqq7u7u7u7vMzMzMzMyZmZl3d3dVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVmZmZVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZVVVVVVVVmZmZVVVVmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3eIiIh3d3dmZmZ3d3d3d3dmZmZ3d3d3d3eIiIiZmZm7u7vMzMzMzMzd3d3d3d3d3d3d3d3MzMzMzMzd3d3d3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3dzMzM3d3d7u7u////////7u7u////////////7u7u////////////////////////////////////////////////////////////////////7u7u3d3d3d3d3d3d3d3d3d3d3d3d3d3dzMzM3d3dzMzM3d3d3d3du7u7u7u7u7u7u7u7qqqqqqqqzMzMzMzMzMzMzMzMu7u7zMzMzMzMzMzM3d3dzMzMzMzMu7u7zMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMzMu7u7u7u7qqqqmZmZmZmZqqqqqqqqqqqqmZmZmZmZqqqqqqqqqqqqqqqqmZmZd3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmd3d3iIiIzMzMzMzMzMzMu7u7zMzMzMzM3d3dqqqqiIiIZmZmZmZmZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmVVVVVVVVVVVVVVVVREREVVVVVVVVZmZmZmZmZmZmd3d3d3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmd3d3ZmZmd3d3iIiImZmZqqqqzMzMzMzM3d3d3d3dzMzM3d3dzMzMzMzM3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7t3d3czMzMzMzO7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///+7u7v///+7u7v///////+7u7t3d3czMzMzMzLu7u8zMzMzMzMzMzMzMzMzMzMzMzN3d3d3d3d3d3e7u7t3d3d3d3d3d3czMzMzMzN3d3d3d3d3d3d3d3d3d3czMzMzMzLu7u8zMzLu7u7u7u6qqqru7u6qqqqqqqqqqqqqqqqqqqqqqqqqqqpmZmYiIiIiIiHd3d3d3d2ZmZmZmZnd3d2ZmZnd3d2ZmZnd3d2ZmZmZmZnd3d4iIiLu7u7u7u8zMzMzMzMzMzLu7u4iIiGZmZmZmZmZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZlVVVWZmZnd3d3d3d4iIiIiIiKqqqqqqqru7u8zMzMzMzMzMzN3d3czMzMzMzN3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////d3d3MzMy7u7vMzMzu7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7MzMzd3d3d3d3d3d3MzMzd3d3d3d3d3d3u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3MzMzd3d3MzMzd3d3MzMzMzMzMzMy7u7u7u7u7u7uqqqqZmZmZmZmZmZl3d3d3d3eIiIiIiIiZmZmIiIiIiIh3d3d3d3d3d3dmZmZmZmZ3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3eIiIiqqqqqqqqqqqqIiIh3d3dmZmZmZmZVVVVVVVVVVVVVVVVERERVVVVVVVVVVVVmZmZVVVVVVVVmZmZmZmZVVVVVVVVVVVVVVVVmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZ3d3eIiIiqqqq7u7u7u7vMzMzMzMzMzMzd3d3MzMzd3d3d3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7uzMzMu7u7u7u73d3d7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u3d3d3d3dzMzMzMzMzMzMzMzM3d3dzMzMzMzMzMzM3d3dzMzMu7u7u7u7u7u7qqqqqqqqmZmZmZmZiIiId3d3d3d3ZmZmZmZmd3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiIiIiId3d3iIiIiIiId3d3iIiId3d3d3d3d3d3d3d3d3d3d3d3ZmZmVVVVVVVVVVVVREREVVVVREREREREVVVVVVVVVVVVVVVVVVVVZmZmVVVVVVVVREREVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVZmZmVVVVZmZmVVVVZmZmVVVVZmZmZmZmZmZmZmZmd3d3mZmZmZmZu7u7zMzMzMzMzMzMzMzMzMzMzMzMzMzM3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD//wAA////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////7u7u3d3du7u7qqqqu7u7zMzM7u7u////////////////////7u7u////////////7u7u////////////////////////////////////////////7u7u////////////////////7u7u////7u7u7u7u7u7u7u7u////7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u7u3d3du7u7u7u7zMzMu7u7u7u7u7u7zMzMu7u7u7u7qqqqqqqqmZmZmZmZmZmZmZmZmZmZiIiIiIiId3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3d3iIiIiIiImZmZiIiIiIiImZmZiIiIiIiIiIiIiIiId3d3d3d3d3d3ZmZmZmZmVVVVVVVVVVVVREREREREREREVVVVREREREREVVVVVVVVVVVVREREVVVVREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmVVVVVVVVZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmd3d3iIiImZmZmZmZqqqqu7u7zMzMzMzMzMzMzMzM3d3dzMzM3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////+7u7u7u7v///////+7u7v///////////////////+7u7v///////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7szMzKqqqpmZmaqqqt3d3d3d3e7u7v///////////////////////////////////////////////////////+7u7v///////////////////+7u7u7u7u7u7u7u7u7u7u7u7t3d3d3d3d3d3d3d3e7u7u7u7t3d3d3d3e7u7t3d3d3d3d3d3d3d3d3d3czMzLu7u7u7u7u7u7u7u6qqqru7u6qqqqqqqpmZmaqqqqqqqpmZmZmZmYiIiIiIiJmZmYiIiIiIiHd3d3d3d4iIiIiIiIiIiHd3d3d3d3d3d4iIiIiIiIiIiHd3d4iIiHd3d3d3d3d3d2ZmZlVVVVVVVVVVVVVVVURERFVVVVVVVURERERERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVVVVVVVVVWZmZlVVVWZmZmZmZmZmZmZmZmZmZlVVVWZmZmZmZmZmZmZmZmZmZmZmZnd3d3d3d3d3d4iIiJmZmaqqqru7u8zMzMzMzMzMzMzMzMzMzMzMzN3d3d3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7d3d27u7uqqqqqqqqqqqrMzMzd3d3u7u7////////////////////////////////u7u7////////////////////////u7u7u7u7u7u7u7u7d3d3d3d3d3d3d3d3d3d3d3d3MzMzMzMzd3d3MzMzMzMzMzMzMzMzd3d3MzMzMzMzMzMzMzMzMzMy7u7u7u7u7u7u7u7u7u7u7u7uqqqq7u7uqqqqZmZmqqqqqqqqqqqqqqqqZmZmqqqqZmZmZmZmIiIiIiIiIiIiIiIiIiIiIiIh3d3d3d3dmZmZ3d3d3d3d3d3dmZmZmZmZVVVVVVVVVVVVEREREREREREREREQzMzNERERERERERERERERERERERERERERVVVVERERVVVVVVVVERERVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3eIiIiZmZmqqqq7u7u7u7u7u7u7u7vMzMzMzMzd3d3d3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u3d3du7u7qqqqmZmZqqqqzMzM3d3d////////////////////////////////////////////////////////////7u7u7u7u7u7u7u7u3d3d3d3d3d3d3d3d3d3dzMzMzMzMzMzMu7u7u7u7u7u7zMzMzMzMu7u7u7u7qqqqu7u7u7u7u7u7qqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqqmZmZmZmZqqqqmZmZmZmZqqqqqqqqmZmZmZmZiIiImZmZiIiId3d3ZmZmZmZmZmZmZmZmZmZmVVVVVVVVVVVVVVVVVVVVVVVVREREREREREREREREREREREREREREREREREREVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmiIiImZmZmZmZqqqqu7u7u7u7u7u7zMzMu7u7zMzM3d3d3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////93d3d3d3bu7u5mZmZmZmaqqqszMzN3d3d3d3e7u7u7u7u7u7u7u7v///+7u7u7u7u7u7t3d3e7u7t3d3d3d3d3d3d3d3d3d3d3d3d3d3czMzN3d3czMzN3d3d3d3czMzMzMzMzMzLu7u6qqqqqqqqqqqpmZmYiIiIiIiIiIiIiIiIiIiHd3d3d3d3d3d4iIiIiIiJmZmZmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d3d3d2ZmZmZmZmZmZlVVVVVVVVVVVVVVVVVVVURERFVVVVVVVURERERERERERERERERERERERFVVVVVVVVVVVVVVVVVVVVVVVVVVVWZmZlVVVWZmZlVVVVVVVVVVVWZmZmZmZnd3d3d3d2ZmZnd3d3d3d3d3d3d3d2ZmZmZmZmZmZmZmZmZmZlVVVVVVVWZmZlVVVWZmZmZmZmZmZnd3d3d3d3d3d3d3d5mZmaqqqru7u7u7u7u7u8zMzMzMzMzMzN3d3d3d3e7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7d3d27u7uqqqqqqqqqqqq7u7u7u7vMzMzd3d3MzMzMzMzMzMzMzMzMzMy7u7u7u7vMzMzMzMzMzMzMzMzMzMzMzMzMzMzd3d3d3d3d3d3d3d3MzMzMzMy7u7uqqqqZmZmIiIiIiIh3d3d3d3dmZmZmZmZmZmZmZmZmZmZmZmZ3d3dmZmZ3d3d3d3d3d3d3d3d3d3dmZmZmZmZmZmZmZmZVVVVVVVVVVVVVVVVVVVVERERERERVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVVmZmZVVVVVVVVVVVVmZmZVVVVmZmZVVVVmZmZVVVVmZmZmZmZmZmZmZmZmZmZmZmZ3d3d3d3d3d3d3d3eIiIiIiIh3d3d3d3d3d3eIiIiIiIhmZmZmZmZmZmZmZmZmZmZmZmZVVVVVVVVmZmZmZmZmZmZ3d3eIiIiIiIiZmZmqqqq7u7u7u7vd3d3MzMzMzMzMzMzd3d3d3d3u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////7u7u7u7u3d3dzMzMu7u7u7u7qqqqqqqqqqqqqqqqqqqqmZmZqqqqqqqqqqqqu7u7u7u7u7u73d3dzMzMzMzMzMzM3d3dzMzM3d3dzMzMzMzMu7u7mZmZmZmZmZmZiIiIiIiIiIiId3d3d3d3d3d3d3d3ZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmVVVVZmZmVVVVVVVVREREVVVVREREVVVVREREVVVVREREVVVVVVVVZmZmVVVVVVVVZmZmZmZmZmZmZmZmZmZmZmZmVVVVZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiImZmZiIiIiIiId3d3iIiIiIiImZmZd3d3d3d3ZmZmZmZmZmZmVVVVVVVVVVVVZmZmd3d3iIiIiIiIiIiImZmZu7u7u7u7zMzMzMzM3d3dzMzM3d3d7u7u7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////+7u7u7u7t3d3d3d3czMzLu7u6qqqqqqqpmZmZmZmZmZmaqqqqqqqqqqqru7u7u7u8zMzLu7u7u7u7u7u7u7u7u7u7u7u7u7u6qqqqqqqqqqqqqqqqqqqoiIiIiIiHd3d2ZmZmZmZlVVVVVVVVVVVURERERERERERERERFVVVURERFVVVURERFVVVVVVVVVVVVVVVWZmZmZmZmZmZmZmZnd3d3d3d3d3d3d3d3d3d3d3d3d3d4iIiIiIiJmZmYiIiIiIiJmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmYiIiJmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmZmYiIiJmZmYiIiHd3d3d3d3d3d2ZmZmZmZnd3d2ZmZmZmZnd3d3d3d3d3d4iIiJmZmaqqqqqqqru7u7u7u8zMzMzMzN3d3d3d3e7u7u7u7v///+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////u7u7////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3d3d3MzMyqqqqqqqqZmZmZmZmZmZmZmZmZmZmqqqqqqqqZmZmqqqqZmZmZmZmZmZmqqqq7u7u7u7u7u7u7u7vMzMy7u7uIiIhVVVVVVVVERERERERERERERERERERERERVVVVVVVVVVVVVVVVmZmZmZmZmZmZ3d3d3d3d3d3eIiIiIiIiIiIiZmZmqqqqZmZmqqqq7u7uqqqq7u7u7u7u7u7vMzMzd3d3MzMzd3d3d3d3d3d3u7u7d3d3u7u7d3d3d3d3MzMzd3d3MzMzd3d3d3d3d3d3d3d3MzMzMzMy7u7uqqqqqqqq7u7uqqqqqqqqqqqqZmZmIiIhmZmZ3d3dmZmZ3d3d3d3eIiIiIiIiZmZmZmZmZmZmZmZm7u7u7u7vMzMzMzMzd3d3d3d3u7u7u7u7u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u3d3dzMzMu7u7u7u7qqqqqqqqmZmZmZmZiIiImZmZiIiImZmZmZmZiIiImZmZmZmZmZmZqqqqqqqqqqqqiIiIZmZmVVVVREREREREVVVVVVVVZmZmZmZmZmZmZmZmd3d3d3d3d3d3iIiIiIiImZmZmZmZqqqqqqqqu7u7zMzM3d3d3d3d3d3d3d3d7u7u7u7u7u7u7u7u7u7u7u7u////////////////////////////////////////////////////////////////7u7u7u7u7u7u3d3d3d3d3d3dzMzMzMzMzMzMu7u7u7u7mZmZmZmZiIiIiIiIiIiImZmZmZmZmZmZqqqqqqqqqqqqmZmZu7u7zMzM3d3d3d3d3d3d7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////+7u7u7u7u7u7t3d3czMzLu7u6qqqqqqqpmZmZmZmZmZmYiIiIiIiIiIiIiIiIiIiIiIiIiIiIiIiHd3d2ZmZlVVVWZmZnd3d3d3d4iIiIiIiIiIiJmZmZmZmaqqqqqqqszMzMzMzMzMzN3d3e7u7u7u7u7u7v///+7u7v///////////////////////////////////////////////////////////////////////////////////////+7u7v///////+7u7v///+7u7v///+7u7u7u7t3d3d3d3d3d3czMzMzMzLu7u7u7u7u7u6qqqru7u7u7u7u7u7u7u7u7u8zMzLu7u8zMzMzMzN3d3e7u7u7u7u7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////u7u7u7u7d3d3MzMzMzMy7u7u7u7uqqqqqqqqqqqqqqqqZmZmZmZmZmZmZmZmZmZmZmZmZmZmqqqq7u7u7u7vMzMzMzMzd3d3d3d3u7u7u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////u7u7u7u7u7u7u7u7u7u7u7u7u7u7d3d3u7u7d3d3d3d3u7u7d3d3u7u7u7u7u7u7u7u7u7u7////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u7u7u3d3d3d3d3d3d3d3dzMzMzMzMzMzMzMzMzMzMzMzM3d3d3d3d3d3d7u7u7u7u7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////7u7u////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7////////////////////u7u7///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+7u7v///////////////////////+7u7v///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////8A////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////7u7u////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AP///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////wD////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////u7u7/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////AW4Akf///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////+mC6TfOQqpjAAAAAElFTkSuQmCC" x="0" y="-452" width="1063px" height="452px" transform="scale(0.0009407338 -0.0022123894)"></svg:image></svg:g></svg:g><svg:g transform=""><svg:text transform="matrix(10.9755 0 0 10.98 425.28 645.8604) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_2" font-size="1px" y="0" x="0" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="0.929" x="-34.227" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="2.0875" x="-32.2918 -31.5688 -31.0678 -30.5108 -30.2318 -29.9528 -29.3958 -28.8388 -28.5598 -28.0588 -27.5018 -27.0008 -26.7218 -26.4428 -25.8858 -25.6068 -25.3838 -24.8268 -24.2698 -23.7128 -23.4338 -23.2108 -22.9318 -22.4308 -22.1518 -21.8728 -21.3158 -20.7588 -20.4798 -19.9228 -19.5888 -19.0318 -18.4748 -17.9178 -17.6948 -17.1938 -16.3598 -16.0808" fill="rgb(0,0,0)">Use the key to identify the organism. </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="4.235" x="-32.2918 -31.7348 -30.3571 -29.7451 -29.1881 -28.6311 -28.3522 -27.5182 -26.9612 -26.4042 -26.1252 -25.5682 -25.2893 -25.0663 -24.5653 -24.2864 -23.7294 -23.4504 -23.1715 -22.8925 -22.3355 -21.7785 -21.4996 -21.2206 -20.8866 -20.3296 -19.7726 -19.4992 -19.2203 -18.6633 -18.3843 -18.1054 -17.8264 -17.2694 -16.7124 -16.4335 -15.8765 -15.3195 -14.7625 -14.2055 -13.9321 -13.6532 -13.3853 -13.1063 -12.8273 -12.5483 -12.2693 -11.9903 -11.7113 -11.4323 -11.1533 -10.8743 -10.5953 -10.3163 -10.0373 -9.7583 -9.4793 -9.2003 -8.9213 -8.6423 -8.3633 -8.0843 -7.8053 -7.5263 -7.2473 -6.9683 -6.6893 -6.4103 -6.1313 -5.8523 -5.5733 -5.2943 -5.0153 -4.7363 -4.4573 -4.1783 -3.8993 -3.6203 -3.3413 -3.0623 -2.7833 -2.5043 -2.2253 -1.9463 -1.6673 -1.3883 -1.1093 -0.8303 -0.5513 -0.2723 0.0067 0.2857 0.5647 0.8437 1.1227 1.4017 1.6807 1.9597 2.2387" fill="rgb(0,0,0)">1 The mouth is at the front of the head.  ........................................................ </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="4.235" x="2.2523 2.5313 3.0885 3.6457 3.9247 4.2039 4.7611 5.0401 5.5973" fill="rgb(0,0,0)"> go to 2 </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="6.2077" x="-32.2918 -30.3564 -29.7443 -29.1872 -28.6301 -28.3511 -27.517 -26.9599 -26.4028 -26.1237 -25.5666 -25.2876 -25.0645 -24.5634 -24.2844 -23.7273 -23.1702 -22.8911 -22.168 -21.6109 -21.0538 -20.4967 -20.2177 -19.9386 -19.3815 -18.8244 -18.5454 -17.9883 -17.4872 -16.9301 -16.6511 -16.094 -15.5369 -14.9798 -14.7008 -14.4217 -13.8646 -13.3075 -13.0285 -12.7494 -12.5263 -11.9692 -11.4681 -11.189 -10.9155 -10.8716 -10.5925 -10.3134 -10.0343 -9.7552 -9.4761 -9.197 -8.9179 -8.6388 -8.3597 -8.0806 -7.8015 -7.5224 -7.2433 -6.9642 -6.6851 -6.406 -6.1269 -5.8478 -5.5687 -5.2896 -5.0105 -4.7314 -4.4523 -4.1732 -3.8941 -3.615 -3.3359 -3.0568 -2.7777 -2.4986 -2.2195 -1.9404 -1.6613 -1.3822 -1.1031 -0.824 -0.5449 -0.2658 0.0133 0.2924 0.5715 0.8506 1.1297 1.4088 1.6879 1.967 2.2461" fill="rgb(0,0,0)"> The mouth is between the eye and the fins.  ............................................... </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="6.2077" x="2.2523" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_3" font-size="1px" y="6.2077" x="2.5311" fill="rgb(0,0,0)">A</svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="6.2077" x="3.2527" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="8.1804" x="-32.2918 -31.7345 -30.3567 -29.7444 -29.1871 -28.6298 -28.3508 -28.1275 -27.5702 -27.0129 -26.4556 -26.1766 -25.8973 -25.674 -25.1167 -24.8432 -24.2859 -23.7286 -23.4496 -23.1703 -22.613 -22.0557 -21.7767 -21.2194 -20.6621 -20.1608 -19.6595 -19.386 -18.8287 -18.2714 -17.7701 -17.4911 -16.9338 -16.3765 -16.1532 -15.5959 -15.3169 -14.8156 -14.2636 -13.7063 -13.427 -12.9257 -12.6464 -12.3729 -12.2743 -11.995 -11.7157 -11.4364 -11.1571 -10.8778 -10.5985 -10.3192 -10.0399 -9.7606 -9.4813 -9.202 -8.9227 -8.6434 -8.3641 -8.0848 -7.8055 -7.5262 -7.2469 -6.9676 -6.6883 -6.409 -6.1297 -5.8504 -5.5711 -5.2918 -5.0125 -4.7332 -4.4539 -4.1746 -3.8953 -3.616 -3.3367 -3.0574 -2.7781 -2.4988 -2.2195 -1.9402 -1.6609 -1.3816 -1.1023 -0.823 -0.5437 -0.2644 0.0149 0.2942 0.5735 0.8528 1.1321 1.4114 1.6907 1.97 2.2493" fill="rgb(0,0,0)">2 The long fin on the back has pale spots.  .................................................... </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="8.1804" x="2.2523 2.5314 3.0887 3.646 3.9251 4.2044 4.7617 5.0408 5.5981" fill="rgb(0,0,0)"> go to 3 </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="10.1531" x="-32.2918 -30.3563 -29.744 -29.1867 -28.6294 -28.2951 -27.7378 -27.4587 -26.9014 -26.5671 -26.0098 -25.7307 -25.1734 -24.6161 -24.337 -23.8357 -23.2784 -22.7211 -22.4418 -21.9405 -21.6614 -21.1041 -20.5468 -20.2677 -19.9941 -19.4365 -18.8792 -18.6001 -18.3768 -17.8195 -17.2622 -16.7049 -16.4258 -16.1465 -15.9232 -15.3659 -15.0866 -14.813 -14.7745 -14.4952 -14.2159 -13.9366 -13.6573 -13.378 -13.0987 -12.8194 -12.5401 -12.2608 -11.9815 -11.7022 -11.4229 -11.1436 -10.8643 -10.585 -10.3057 -10.0264 -9.7471 -9.4678 -9.1885 -8.9092 -8.6299 -8.3506 -8.0713 -7.792 -7.5127 -7.2334 -6.9541 -6.6748 -6.3955 -6.1162 -5.8369 -5.5576 -5.2783 -4.999 -4.7197 -4.4404 -4.1611 -3.8818 -3.6025 -3.3232 -3.0439 -2.7646 -2.4853 -2.206 -1.9267 -1.6474 -1.3681 -1.0888 -0.8095 -0.5302 -0.2509 0.0284 0.3077 0.587 0.8663 1.1456 1.4249 1.7042 1.9835 2.2628" fill="rgb(0,0,0)"> There are no spots on the long fin.  ............................................................. </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="10.1531" x="2.2523" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_3" font-size="1px" y="10.1531" x="2.5311" fill="rgb(0,0,0)">B</svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="10.1531" x="3.2527" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="12.1203" x="-32.2918 -31.7347 -30.3569 -29.7448 -29.1877 -28.6306 -28.3516 -28.0725 -27.5154 -27.2923 -27.0692 -26.7902 -26.5111 -26.288 -25.7309 -25.4574 -25.2343 -24.7332 -24.4542 -24.2311 -23.674 -23.1169 -22.5598 -22.0027 -21.6686 -21.3896 -21.1105 -20.5534 -20.0014 -19.4439 -19.1649 -18.8858 -18.3287 -17.7716 -17.4926 -16.9355 -16.3784 -15.8213 -15.3202 -15.0411 -14.7621 -14.4941 -14.215 -13.9359 -13.6568 -13.3777 -13.0986 -12.8195 -12.5404 -12.2613 -11.9822 -11.7031 -11.424 -11.1449 -10.8658 -10.5867 -10.3076 -10.0285 -9.7494 -9.4703 -9.1912 -8.9121 -8.633 -8.3539 -8.0748 -7.7957 -7.5166 -7.2375 -6.9584 -6.6793 -6.4002 -6.1211 -5.842 -5.5629 -5.2838 -5.0047 -4.7256 -4.4465 -4.1674 -3.8883 -3.6092 -3.3301 -3.051 -2.7719 -2.4928 -2.2137 -1.9346 -1.6555 -1.3764 -1.0973 -0.8182 -0.5391 -0.26 0.0191 0.2982 0.5773 0.8564 1.1355 1.4146 1.6937 1.9728 2.2519" fill="rgb(0,0,0)">3 The tail fin is longer than the body.  ............................................................ </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="12.1203" x="2.2523" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_3" font-size="1px" y="12.1203" x="2.5311" fill="rgb(0,0,0)">C</svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="12.1203" x="3.2527" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="14.093" x="-32.2918 -30.351 -29.7389 -29.1818 -28.6247 -28.3457 -28.0666 -27.5095 -27.2864 -27.0633 -26.7843 -26.5052 -26.2821 -25.725 -25.4515 -25.2284 -24.7273 -24.4483 -23.9472 -23.3901 -22.833 -22.4989 -22.2198 -21.6627 -21.3286 -21.0496 -20.7705 -20.2134 -19.6614 -19.1039 -18.8249 -18.5458 -17.9887 -17.4316 -17.1526 -16.5955 -16.0384 -15.4813 -14.9802 -14.7011 -14.4221 -14.2142 -13.9351 -13.656 -13.3769 -13.0978 -12.8187 -12.5396 -12.2605 -11.9814 -11.7023 -11.4232 -11.1441 -10.865 -10.5859 -10.3068 -10.0277 -9.7486 -9.4695 -9.1904 -8.9113 -8.6322 -8.3531 -8.074 -7.7949 -7.5158 -7.2367 -6.9576 -6.6785 -6.3994 -6.1203 -5.8412 -5.5621 -5.283 -5.0039 -4.7248 -4.4457 -4.1666 -3.8875 -3.6084 -3.3293 -3.0502 -2.7711 -2.492 -2.2129 -1.9338 -1.6547 -1.3756 -1.0965 -0.8174 -0.5383 -0.2592 0.0199 0.299 0.5781 0.8572 1.1363 1.4154 1.6945 1.9736 2.2527" fill="rgb(0,0,0)"> The tail fin is shorter than the body.  ........................................................... </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="14.093" x="2.2523" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_3" font-size="1px" y="14.093" x="2.5311" fill="rgb(0,0,0)">D</svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="14.093" x="3.2527" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="15.246" x="-34.227" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="16.399" x="-34.227" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_3" font-size="1px" y="17.552" x="-34.227" fill="rgb(0,0,0)">4</svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="17.552" x="-33.6694 -32.2916 -31.3462 -30.7888 -30.5654 -30.064 -29.5066 -29.2276 -28.9482 -28.3908 -27.8334 -27.554 -27.002 -26.6685 -26.1111 -25.6097 -25.3307 -24.7733 -24.4389 -23.8815 -23.6025 -23.0451 -22.4877 -21.9863 -21.4849 -20.9275 -20.4261 -19.9247 -19.3673 -18.8099 -18.5309 -17.9735 -17.4721" fill="rgb(0,0,0)"> Which features are possessed by </svg:tspan><svg:tspan font-family="g_font_3" font-size="1px" y="17.552" x="-17.1928 -16.6356 -16.3564" fill="rgb(0,0,0)">all</svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="17.552" x="-16.0776 -15.7986 -15.2408 -15.017 -14.4592 -13.9014 -13.6216 -13.3426 -12.8408 -12.283 -12.0645 -11.8405 -11.3387 -10.7867" fill="rgb(0,0,0)"> plant cells? </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="18.6995" x="-34.227" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="20.2022" x="-30.9962 -28.4048 -27.8471 -27.5681 -27.0664 -26.5087 -26.285 -26.0613 -25.7823 -25.0586 -24.5009 -24.2772 -24.0587 -21.9593 -21.4576 -20.8999 -20.6762 -20.1185 -19.7838 -19.2261 -18.6684 -18.4447 -17.887 -17.3853 -17.1118 -16.6143" fill="rgb(0,0,0)"> a cell wall chloroplasts </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="19.9017" x="-12.3384" fill="rgb(0,0,0)"> </svg:tspan></svg:text></svg:g><svg:g transform=""><svg:path d="M 70.68 438.08 L 71.16 438.08 L 71.16 437.6 L 70.68 437.6 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 70.68 438.08 L 252 438.08 L 252 437.6 L 70.68 437.6 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 251.52 438.08 L 252 438.08 L 252 437.6 L 251.52 437.6 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 70.68 437.6 L 71.16 437.6 L 71.16 418.22 L 70.68 418.22 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 99.06 437.6 L 99.54 437.6 L 99.54 418.22 L 99.06 418.22 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 175.26 437.6 L 175.74 437.6 L 175.74 418.22 L 175.26 418.22 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 251.52 437.6 L 252 437.6 L 252 418.22 L 251.52 418.22 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:text transform="matrix(10.9755 0 0 10.98 81.12 400.9403) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_3" font-size="1px" y="0" x="0 0.7214" fill="rgb(0,0,0)">A </svg:tspan><svg:tspan font-family="g_font_8" font-size="1px" y="0" x="4.6686" fill="rgb(0,0,0)"></svg:tspan><svg:tspan font-family="g_font_9" font-size="1px" y="0" x="5.5815" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_8" font-size="1px" y="0" x="11.6167" fill="rgb(0,0,0)"></svg:tspan><svg:tspan font-family="g_font_9" font-size="1px" y="0" x="12.5296" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="0" x="16.0392 16.5414 17.0996 17.5971" fill="rgb(0,0,0)">key </svg:tspan></svg:text></svg:g><svg:g transform=""><svg:path d="M 70.68 418.22 L 252 418.22 L 252 417.74 L 70.68 417.74 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 70.68 417.74 L 71.16 417.74 L 71.16 396.74 L 70.68 396.74 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 99.06 417.74 L 99.54 417.74 L 99.54 396.74 L 99.06 396.74 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 175.26 417.74 L 175.74 417.74 L 175.74 396.74 L 175.26 396.74 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 251.52 417.74 L 252 417.74 L 252 396.74 L 251.52 396.74 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:text transform="matrix(10.9755 0 0 10.98 81.12 379.9403) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_3" font-size="1px" y="0" x="0 0.7214" fill="rgb(0,0,0)">B </svg:tspan><svg:tspan font-family="g_font_8" font-size="1px" y="0" x="4.6686" fill="rgb(0,0,0)"></svg:tspan><svg:tspan font-family="g_font_9" font-size="1px" y="0" x="5.5815" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_8" font-size="1px" y="0" x="11.6167" fill="rgb(0,0,0)"></svg:tspan><svg:tspan font-family="g_font_9" font-size="1px" y="0" x="12.5296" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_8" font-size="1px" y="0" x="16.0392" fill="rgb(0,0,0)"></svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="0" x="16.9521 17.5374 17.8164 18.3737 18.708 19.2653 19.7666 20.3239 20.8812 21.1605" fill="rgb(0,0,0)">= present </svg:tspan></svg:text></svg:g><svg:g transform=""><svg:path d="M 70.68 396.74 L 71.16 396.74 L 71.16 375.74 L 70.68 375.74 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 99.06 396.74 L 99.54 396.74 L 99.54 375.74 L 99.06 375.74 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 175.26 396.74 L 175.74 396.74 L 175.74 375.74 L 175.26 375.74 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 251.52 396.74 L 252 396.74 L 252 375.74 L 251.52 375.74 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:text transform="matrix(10.9755 0 0 10.98 81.12 358.9403) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_3" font-size="1px" y="0" x="0 0.7214" fill="rgb(0,0,0)">C </svg:tspan><svg:tspan font-family="g_font_8" font-size="1px" y="0" x="4.6686" fill="rgb(0,0,0)"></svg:tspan><svg:tspan font-family="g_font_9" font-size="1px" y="0" x="5.5815" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_8" font-size="1px" y="0" x="11.6167" fill="rgb(0,0,0)"></svg:tspan><svg:tspan font-family="g_font_9" font-size="1px" y="0" x="12.5296" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_8" font-size="1px" y="0" x="16.0392" fill="rgb(0,0,0)"></svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="0" x="16.9521 17.5376 17.8166 18.3741 18.9316 19.4331 19.9906 20.5481 20.8216" fill="rgb(0,0,0)">= absent </svg:tspan></svg:text></svg:g><svg:g transform=""><svg:path d="M 70.68 375.74 L 71.16 375.74 L 71.16 354.74 L 70.68 354.74 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 99.06 375.74 L 99.54 375.74 L 99.54 354.74 L 99.06 354.74 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 175.26 375.74 L 175.74 375.74 L 175.74 354.74 L 175.26 354.74 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 251.52 375.74 L 252 375.74 L 252 354.74 L 251.52 354.74 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:text transform="matrix(10.9755 0 0 10.98 81.12 337.9403) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_3" font-size="1px" y="0" x="0 0.7214" fill="rgb(0,0,0)">D </svg:tspan><svg:tspan font-family="g_font_8" font-size="1px" y="0" x="4.6686" fill="rgb(0,0,0)"></svg:tspan><svg:tspan font-family="g_font_9" font-size="1px" y="0" x="5.5815" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_8" font-size="1px" y="0" x="11.6167" fill="rgb(0,0,0)"></svg:tspan><svg:tspan font-family="g_font_9" font-size="1px" y="0" x="12.5296 16.0394" fill="rgb(0,0,0)">  </svg:tspan></svg:text></svg:g><svg:g transform=""><svg:path d="M 70.68 354.74 L 71.16 354.74 L 71.16 333.2 L 70.68 333.2 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 70.68 333.68 L 99.06 333.68 L 99.06 333.2 L 70.68 333.2 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 99.06 354.74 L 99.54 354.74 L 99.54 333.2 L 99.06 333.2 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 99.54 333.68 L 175.26 333.68 L 175.26 333.2 L 99.54 333.2 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 175.26 354.74 L 175.74 354.74 L 175.74 333.2 L 175.26 333.2 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 175.74 333.68 L 251.52 333.68 L 251.52 333.2 L 175.74 333.2 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 251.52 354.74 L 252 354.74 L 252 333.2 L 251.52 333.2 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:path d="M 251.52 333.68 L 252 333.68 L 252 333.2 L 251.52 333.2 Z" stroke-miterlimit="0" stroke-linecap="" stroke-linejoin="" stroke-width="1px" stroke-dasharray="" stroke-dashoffset="0px" fill="rgb(0,0,0)"></svg:path><svg:text transform="matrix(10.9755 0 0 10.98 49.62 323.0004) scale(1, -1)" xml:space="preserve"><svg:tspan font-family="g_font_2" font-size="1px" y="0" x="0" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="1.153" x="0" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_3" font-size="1px" y="2.306" x="0" fill="rgb(0,0,0)">5</svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="2.306" x="0.5576 1.9354 2.8808 3.4382 3.6616 4.163 4.7204 4.9994 5.2228 5.7802 6.2816 6.839 7.0624 7.3359 7.8933 8.1727 8.4517 9.0091 9.3435 9.9009 10.4583 11.0157 11.2391 11.7405 12.2979 12.5773 12.8007 13.3581 13.9155 14.1945 14.4179 14.9193 15.1983 15.6997 16.2571 16.8145 17.5379 18.0953 18.3688 18.9262 19.4276 19.7066 19.986 20.5434 21.1008 21.3798 21.9372 22.4946 22.996 23.5534 24.1108 24.6682 25.2256 25.783 26.3404 26.8418 27.1212 27.4002 27.9576 28.515 29.067 29.5699 29.9043 30.4617 31.0191 31.5205 31.7999 32.0789 32.5803 32.8597 33.4171 34.2426 34.8 35.3014 35.8588 36.1378 36.6952 37.2526 37.81 38.089 38.3124 38.5358 39.0372 39.5892 39.9227 40.4801" fill="rgb(0,0,0)"> Which level of organisation is shown by the oesophagus, pancreas, stomach and liver? </svg:tspan><svg:tspan font-family="g_font_3" font-size="1px" y="4.459" x="1.9352 2.6566" fill="rgb(0,0,0)">A </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="4.459" x="3.8704 4.3716 4.9288 5.152 5.3752 5.8764" fill="rgb(0,0,0)">cells </svg:tspan><svg:tspan font-family="g_font_3" font-size="1px" y="6.4262" x="1.9352 2.6566" fill="rgb(0,0,0)">B </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="6.4262" x="3.8704 4.428 4.7626 5.3202 5.8778 6.4354 6.937" fill="rgb(0,0,0)">organs </svg:tspan><svg:tspan font-family="g_font_3" font-size="1px" y="8.3989" x="1.9352 2.6566" fill="rgb(0,0,0)">C </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="8.3989" x="3.8704 4.4279 4.7624 5.3199 5.8774 6.4349 6.6584 7.1599 7.9944 8.4959" fill="rgb(0,0,0)">organisms </svg:tspan><svg:tspan font-family="g_font_3" font-size="1px" y="10.3716" x="1.9407 2.6621" fill="rgb(0,0,0)">D </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="10.3716" x="3.8759 4.1558 4.3797 4.8816 5.3835 5.9414 6.4993 6.9968" fill="rgb(0,0,0)">tissues </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="11.5246" x="0" fill="rgb(0,0,0)"> </svg:tspan><svg:tspan font-family="g_font_2" font-size="1px" y="12.6776" x="0" fill="rgb(0,0,0)"> </svg:tspan></svg:text></svg:g></svg:g></svg:svg>